module PLIC(
  input   clk,
  input   reset,
  input   io_devices_0_valid,
  output  io_devices_0_ready,
  output  io_devices_0_complete,
  input   io_devices_1_valid,
  output  io_devices_1_ready,
  output  io_devices_1_complete,
  input   io_devices_2_valid,
  output  io_devices_2_ready,
  output  io_devices_2_complete,
  input   io_devices_3_valid,
  output  io_devices_3_ready,
  output  io_devices_3_complete,
  input   io_devices_4_valid,
  output  io_devices_4_ready,
  output  io_devices_4_complete,
  input   io_devices_5_valid,
  output  io_devices_5_ready,
  output  io_devices_5_complete,
  input   io_devices_6_valid,
  output  io_devices_6_ready,
  output  io_devices_6_complete,
  input   io_devices_7_valid,
  output  io_devices_7_ready,
  output  io_devices_7_complete,
  input   io_devices_8_valid,
  output  io_devices_8_ready,
  output  io_devices_8_complete,
  input   io_devices_9_valid,
  output  io_devices_9_ready,
  output  io_devices_9_complete,
  input   io_devices_10_valid,
  output  io_devices_10_ready,
  output  io_devices_10_complete,
  input   io_devices_11_valid,
  output  io_devices_11_ready,
  output  io_devices_11_complete,
  input   io_devices_12_valid,
  output  io_devices_12_ready,
  output  io_devices_12_complete,
  input   io_devices_13_valid,
  output  io_devices_13_ready,
  output  io_devices_13_complete,
  input   io_devices_14_valid,
  output  io_devices_14_ready,
  output  io_devices_14_complete,
  input   io_devices_15_valid,
  output  io_devices_15_ready,
  output  io_devices_15_complete,
  input   io_devices_16_valid,
  output  io_devices_16_ready,
  output  io_devices_16_complete,
  input   io_devices_17_valid,
  output  io_devices_17_ready,
  output  io_devices_17_complete,
  input   io_devices_18_valid,
  output  io_devices_18_ready,
  output  io_devices_18_complete,
  input   io_devices_19_valid,
  output  io_devices_19_ready,
  output  io_devices_19_complete,
  input   io_devices_20_valid,
  output  io_devices_20_ready,
  output  io_devices_20_complete,
  input   io_devices_21_valid,
  output  io_devices_21_ready,
  output  io_devices_21_complete,
  input   io_devices_22_valid,
  output  io_devices_22_ready,
  output  io_devices_22_complete,
  input   io_devices_23_valid,
  output  io_devices_23_ready,
  output  io_devices_23_complete,
  input   io_devices_24_valid,
  output  io_devices_24_ready,
  output  io_devices_24_complete,
  input   io_devices_25_valid,
  output  io_devices_25_ready,
  output  io_devices_25_complete,
  input   io_devices_26_valid,
  output  io_devices_26_ready,
  output  io_devices_26_complete,
  input   io_devices_27_valid,
  output  io_devices_27_ready,
  output  io_devices_27_complete,
  input   io_devices_28_valid,
  output  io_devices_28_ready,
  output  io_devices_28_complete,
  input   io_devices_29_valid,
  output  io_devices_29_ready,
  output  io_devices_29_complete,
  input   io_devices_30_valid,
  output  io_devices_30_ready,
  output  io_devices_30_complete,
  output  io_harts_0,
  output  io_tl_acquire_ready,
  input   io_tl_acquire_valid,
  input  [25:0] io_tl_acquire_bits_addr_block,
  input  [1:0] io_tl_acquire_bits_client_xact_id,
  input  [2:0] io_tl_acquire_bits_addr_beat,
  input   io_tl_acquire_bits_is_builtin_type,
  input  [2:0] io_tl_acquire_bits_a_type,
  input  [11:0] io_tl_acquire_bits_union,
  input  [63:0] io_tl_acquire_bits_data,
  input   io_tl_grant_ready,
  output  io_tl_grant_valid,
  output [2:0] io_tl_grant_bits_addr_beat,
  output [1:0] io_tl_grant_bits_client_xact_id,
  output  io_tl_grant_bits_manager_xact_id,
  output  io_tl_grant_bits_is_builtin_type,
  output [3:0] io_tl_grant_bits_g_type,
  output [63:0] io_tl_grant_bits_data
);
  wire  T_680_0;
  wire  T_680_1;
  wire  T_680_2;
  wire  T_680_3;
  wire  T_680_4;
  wire  T_680_5;
  wire  T_680_6;
  wire  T_680_7;
  wire  T_680_8;
  wire  T_680_9;
  wire  T_680_10;
  wire  T_680_11;
  wire  T_680_12;
  wire  T_680_13;
  wire  T_680_14;
  wire  T_680_15;
  wire  T_680_16;
  wire  T_680_17;
  wire  T_680_18;
  wire  T_680_19;
  wire  T_680_20;
  wire  T_680_21;
  wire  T_680_22;
  wire  T_680_23;
  wire  T_680_24;
  wire  T_680_25;
  wire  T_680_26;
  wire  T_680_27;
  wire  T_680_28;
  wire  T_680_29;
  wire  T_680_30;
  wire  T_680_31;
  wire  priority_0;
  wire  priority_1;
  wire  priority_2;
  wire  priority_3;
  wire  priority_4;
  wire  priority_5;
  wire  priority_6;
  wire  priority_7;
  wire  priority_8;
  wire  priority_9;
  wire  priority_10;
  wire  priority_11;
  wire  priority_12;
  wire  priority_13;
  wire  priority_14;
  wire  priority_15;
  wire  priority_16;
  wire  priority_17;
  wire  priority_18;
  wire  priority_19;
  wire  priority_20;
  wire  priority_21;
  wire  priority_22;
  wire  priority_23;
  wire  priority_24;
  wire  priority_25;
  wire  priority_26;
  wire  priority_27;
  wire  priority_28;
  wire  priority_29;
  wire  priority_30;
  wire  priority_31;
  wire  T_691_0;
  wire  threshold_0;
  wire  T_733_0;
  wire  T_733_1;
  wire  T_733_2;
  wire  T_733_3;
  wire  T_733_4;
  wire  T_733_5;
  wire  T_733_6;
  wire  T_733_7;
  wire  T_733_8;
  wire  T_733_9;
  wire  T_733_10;
  wire  T_733_11;
  wire  T_733_12;
  wire  T_733_13;
  wire  T_733_14;
  wire  T_733_15;
  wire  T_733_16;
  wire  T_733_17;
  wire  T_733_18;
  wire  T_733_19;
  wire  T_733_20;
  wire  T_733_21;
  wire  T_733_22;
  wire  T_733_23;
  wire  T_733_24;
  wire  T_733_25;
  wire  T_733_26;
  wire  T_733_27;
  wire  T_733_28;
  wire  T_733_29;
  wire  T_733_30;
  wire  T_733_31;
  reg  pending_0;
  reg [31:0] GEN_100;
  reg  pending_1;
  reg [31:0] GEN_132;
  reg  pending_2;
  reg [31:0] GEN_133;
  reg  pending_3;
  reg [31:0] GEN_227;
  reg  pending_4;
  reg [31:0] GEN_259;
  reg  pending_5;
  reg [31:0] GEN_260;
  reg  pending_6;
  reg [31:0] GEN_292;
  reg  pending_7;
  reg [31:0] GEN_293;
  reg  pending_8;
  reg [31:0] GEN_325;
  reg  pending_9;
  reg [31:0] GEN_327;
  reg  pending_10;
  reg [31:0] GEN_328;
  reg  pending_11;
  reg [31:0] GEN_360;
  reg  pending_12;
  reg [31:0] GEN_361;
  reg  pending_13;
  reg [31:0] GEN_393;
  reg  pending_14;
  reg [31:0] GEN_394;
  reg  pending_15;
  reg [31:0] GEN_395;
  reg  pending_16;
  reg [31:0] GEN_396;
  reg  pending_17;
  reg [31:0] GEN_397;
  reg  pending_18;
  reg [31:0] GEN_399;
  reg  pending_19;
  reg [31:0] GEN_400;
  reg  pending_20;
  reg [31:0] GEN_402;
  reg  pending_21;
  reg [31:0] GEN_403;
  reg  pending_22;
  reg [31:0] GEN_405;
  reg  pending_23;
  reg [31:0] GEN_406;
  reg  pending_24;
  reg [31:0] GEN_408;
  reg  pending_25;
  reg [31:0] GEN_409;
  reg  pending_26;
  reg [31:0] GEN_411;
  reg  pending_27;
  reg [31:0] GEN_412;
  reg  pending_28;
  reg [31:0] GEN_414;
  reg  pending_29;
  reg [31:0] GEN_415;
  reg  pending_30;
  reg [31:0] GEN_417;
  reg  pending_31;
  reg [31:0] GEN_418;
  reg  enables_0_0;
  reg [31:0] GEN_420;
  reg  enables_0_1;
  reg [31:0] GEN_421;
  reg  enables_0_2;
  reg [31:0] GEN_423;
  reg  enables_0_3;
  reg [31:0] GEN_424;
  reg  enables_0_4;
  reg [31:0] GEN_426;
  reg  enables_0_5;
  reg [31:0] GEN_427;
  reg  enables_0_6;
  reg [31:0] GEN_429;
  reg  enables_0_7;
  reg [31:0] GEN_430;
  reg  enables_0_8;
  reg [31:0] GEN_432;
  reg  enables_0_9;
  reg [31:0] GEN_433;
  reg  enables_0_10;
  reg [31:0] GEN_435;
  reg  enables_0_11;
  reg [31:0] GEN_436;
  reg  enables_0_12;
  reg [31:0] GEN_438;
  reg  enables_0_13;
  reg [31:0] GEN_439;
  reg  enables_0_14;
  reg [31:0] GEN_441;
  reg  enables_0_15;
  reg [31:0] GEN_442;
  reg  enables_0_16;
  reg [31:0] GEN_444;
  reg  enables_0_17;
  reg [31:0] GEN_445;
  reg  enables_0_18;
  reg [31:0] GEN_447;
  reg  enables_0_19;
  reg [31:0] GEN_448;
  reg  enables_0_20;
  reg [31:0] GEN_450;
  reg  enables_0_21;
  reg [31:0] GEN_451;
  reg  enables_0_22;
  reg [31:0] GEN_453;
  reg  enables_0_23;
  reg [31:0] GEN_454;
  reg  enables_0_24;
  reg [31:0] GEN_456;
  reg  enables_0_25;
  reg [31:0] GEN_457;
  reg  enables_0_26;
  reg [31:0] GEN_459;
  reg  enables_0_27;
  reg [31:0] GEN_460;
  reg  enables_0_28;
  reg [31:0] GEN_462;
  reg  enables_0_29;
  reg [31:0] GEN_463;
  reg  enables_0_30;
  reg [31:0] GEN_465;
  reg  enables_0_31;
  reg [31:0] GEN_466;
  wire  T_770;
  wire  GEN_69;
  wire  T_774;
  wire  GEN_70;
  wire  T_778;
  wire  GEN_71;
  wire  T_782;
  wire  GEN_72;
  wire  T_786;
  wire  GEN_73;
  wire  T_790;
  wire  GEN_74;
  wire  T_794;
  wire  GEN_75;
  wire  T_798;
  wire  GEN_76;
  wire  T_802;
  wire  GEN_77;
  wire  T_806;
  wire  GEN_78;
  wire  T_810;
  wire  GEN_79;
  wire  T_814;
  wire  GEN_80;
  wire  T_818;
  wire  GEN_81;
  wire  T_822;
  wire  GEN_82;
  wire  T_826;
  wire  GEN_83;
  wire  T_830;
  wire  GEN_84;
  wire  T_834;
  wire  GEN_85;
  wire  T_838;
  wire  GEN_86;
  wire  T_842;
  wire  GEN_87;
  wire  T_846;
  wire  GEN_88;
  wire  T_850;
  wire  GEN_89;
  wire  T_854;
  wire  GEN_90;
  wire  T_858;
  wire  GEN_91;
  wire  T_862;
  wire  GEN_92;
  wire  T_866;
  wire  GEN_93;
  wire  T_870;
  wire  GEN_94;
  wire  T_874;
  wire  GEN_95;
  wire  T_878;
  wire  GEN_96;
  wire  T_882;
  wire  GEN_97;
  wire  T_886;
  wire  GEN_98;
  wire  T_890;
  wire  GEN_99;
  wire [4:0] maxDevs_0;
  wire  T_900;
  wire [1:0] T_901;
  wire  T_902;
  wire [1:0] T_903;
  wire  T_904;
  wire [1:0] T_905;
  wire  T_906;
  wire [1:0] T_907;
  wire  T_908;
  wire [1:0] T_909;
  wire  T_910;
  wire [1:0] T_911;
  wire  T_912;
  wire [1:0] T_913;
  wire  T_914;
  wire [1:0] T_915;
  wire  T_916;
  wire [1:0] T_917;
  wire  T_918;
  wire [1:0] T_919;
  wire  T_920;
  wire [1:0] T_921;
  wire  T_922;
  wire [1:0] T_923;
  wire  T_924;
  wire [1:0] T_925;
  wire  T_926;
  wire [1:0] T_927;
  wire  T_928;
  wire [1:0] T_929;
  wire  T_930;
  wire [1:0] T_931;
  wire  T_932;
  wire [1:0] T_933;
  wire  T_934;
  wire [1:0] T_935;
  wire  T_936;
  wire [1:0] T_937;
  wire  T_938;
  wire [1:0] T_939;
  wire  T_940;
  wire [1:0] T_941;
  wire  T_942;
  wire [1:0] T_943;
  wire  T_944;
  wire [1:0] T_945;
  wire  T_946;
  wire [1:0] T_947;
  wire  T_948;
  wire [1:0] T_949;
  wire  T_950;
  wire [1:0] T_951;
  wire  T_952;
  wire [1:0] T_953;
  wire  T_954;
  wire [1:0] T_955;
  wire  T_956;
  wire [1:0] T_957;
  wire  T_958;
  wire [1:0] T_959;
  wire  T_960;
  wire [1:0] T_961;
  wire  T_966;
  wire [1:0] T_967;
  wire [1:0] T_969;
  wire  T_970;
  wire  T_971;
  wire  T_974;
  wire [1:0] T_975;
  wire  T_979;
  wire  T_980;
  wire [1:0] T_981;
  wire [1:0] GEN_702;
  wire [2:0] T_983;
  wire [1:0] T_984;
  wire [1:0] T_985;
  wire  T_988;
  wire [1:0] T_989;
  wire  T_993;
  wire  T_996;
  wire [1:0] T_997;
  wire  T_1001;
  wire  T_1002;
  wire [1:0] T_1003;
  wire [1:0] GEN_703;
  wire [2:0] T_1005;
  wire [1:0] T_1006;
  wire [1:0] T_1007;
  wire  T_1008;
  wire [1:0] T_1009;
  wire [2:0] GEN_704;
  wire [3:0] T_1011;
  wire [2:0] T_1012;
  wire [2:0] T_1013;
  wire  T_1016;
  wire [1:0] T_1017;
  wire  T_1021;
  wire  T_1024;
  wire [1:0] T_1025;
  wire  T_1029;
  wire  T_1030;
  wire [1:0] T_1031;
  wire [1:0] GEN_705;
  wire [2:0] T_1033;
  wire [1:0] T_1034;
  wire [1:0] T_1035;
  wire  T_1038;
  wire [1:0] T_1039;
  wire  T_1043;
  wire  T_1046;
  wire [1:0] T_1047;
  wire  T_1051;
  wire  T_1052;
  wire [1:0] T_1053;
  wire [1:0] GEN_706;
  wire [2:0] T_1055;
  wire [1:0] T_1056;
  wire [1:0] T_1057;
  wire  T_1058;
  wire [1:0] T_1059;
  wire [2:0] GEN_707;
  wire [3:0] T_1061;
  wire [2:0] T_1062;
  wire [2:0] T_1063;
  wire  T_1064;
  wire [1:0] T_1065;
  wire [3:0] GEN_708;
  wire [4:0] T_1067;
  wire [3:0] T_1068;
  wire [3:0] T_1069;
  wire  T_1072;
  wire [1:0] T_1073;
  wire  T_1077;
  wire  T_1080;
  wire [1:0] T_1081;
  wire  T_1085;
  wire  T_1086;
  wire [1:0] T_1087;
  wire [1:0] GEN_709;
  wire [2:0] T_1089;
  wire [1:0] T_1090;
  wire [1:0] T_1091;
  wire  T_1094;
  wire [1:0] T_1095;
  wire  T_1099;
  wire  T_1102;
  wire [1:0] T_1103;
  wire  T_1107;
  wire  T_1108;
  wire [1:0] T_1109;
  wire [1:0] GEN_710;
  wire [2:0] T_1111;
  wire [1:0] T_1112;
  wire [1:0] T_1113;
  wire  T_1114;
  wire [1:0] T_1115;
  wire [2:0] GEN_711;
  wire [3:0] T_1117;
  wire [2:0] T_1118;
  wire [2:0] T_1119;
  wire  T_1122;
  wire [1:0] T_1123;
  wire  T_1127;
  wire  T_1130;
  wire [1:0] T_1131;
  wire  T_1135;
  wire  T_1136;
  wire [1:0] T_1137;
  wire [1:0] GEN_712;
  wire [2:0] T_1139;
  wire [1:0] T_1140;
  wire [1:0] T_1141;
  wire  T_1144;
  wire [1:0] T_1145;
  wire  T_1149;
  wire  T_1152;
  wire [1:0] T_1153;
  wire  T_1157;
  wire  T_1158;
  wire [1:0] T_1159;
  wire [1:0] GEN_713;
  wire [2:0] T_1161;
  wire [1:0] T_1162;
  wire [1:0] T_1163;
  wire  T_1164;
  wire [1:0] T_1165;
  wire [2:0] GEN_714;
  wire [3:0] T_1167;
  wire [2:0] T_1168;
  wire [2:0] T_1169;
  wire  T_1170;
  wire [1:0] T_1171;
  wire [3:0] GEN_715;
  wire [4:0] T_1173;
  wire [3:0] T_1174;
  wire [3:0] T_1175;
  wire  T_1176;
  wire [1:0] T_1177;
  wire [4:0] GEN_716;
  wire [5:0] T_1179;
  wire [4:0] T_1180;
  wire [4:0] T_1181;
  reg [4:0] T_1182;
  reg [31:0] GEN_468;
  reg [1:0] T_1183;
  reg [31:0] GEN_469;
  wire [1:0] T_1185;
  wire  T_1186;
  wire  acq_clk;
  wire  acq_reset;
  wire  acq_io_enq_ready;
  wire  acq_io_enq_valid;
  wire [25:0] acq_io_enq_bits_addr_block;
  wire [1:0] acq_io_enq_bits_client_xact_id;
  wire [2:0] acq_io_enq_bits_addr_beat;
  wire  acq_io_enq_bits_is_builtin_type;
  wire [2:0] acq_io_enq_bits_a_type;
  wire [11:0] acq_io_enq_bits_union;
  wire [63:0] acq_io_enq_bits_data;
  wire  acq_io_deq_ready;
  wire  acq_io_deq_valid;
  wire [25:0] acq_io_deq_bits_addr_block;
  wire [1:0] acq_io_deq_bits_client_xact_id;
  wire [2:0] acq_io_deq_bits_addr_beat;
  wire  acq_io_deq_bits_is_builtin_type;
  wire [2:0] acq_io_deq_bits_a_type;
  wire [11:0] acq_io_deq_bits_union;
  wire [63:0] acq_io_deq_bits_data;
  wire  acq_io_count;
  wire  T_1210;
  wire  T_1212;
  wire  T_1213;
  wire  read;
  wire  T_1216;
  wire  T_1217;
  wire  write;
  wire  T_1220;
  wire  T_1221;
  wire  T_1222;
  wire  T_1223;
  wire  T_1225;
  wire [2:0] T_1233_0;
  wire [2:0] T_1233_1;
  wire  T_1235;
  wire  T_1236;
  wire  T_1237;
  wire  T_1238;
  wire [2:0] T_1239;
  wire [2:0] T_1241;
  wire [28:0] T_1242;
  wire [31:0] T_1243;
  wire [25:0] addr;
  wire  hart;
  wire [4:0] GEN_0;
  wire [5:0] T_1245;
  wire [4:0] myMaxDev;
  wire [63:0] rdata;
  wire  T_1251;
  wire  T_1252;
  wire  T_1254;
  wire [1:0] T_1256;
  wire  T_1257;
  wire  T_1258;
  wire [3:0] T_1262;
  wire [3:0] T_1266;
  wire [7:0] T_1267;
  wire  T_1269;
  wire  T_1270;
  wire  T_1274;
  wire [7:0] T_1275;
  wire [7:0] T_1277;
  wire [7:0] T_1278;
  wire  T_1279;
  wire  T_1280;
  wire  T_1281;
  wire  T_1282;
  wire  T_1283;
  wire  T_1284;
  wire  T_1285;
  wire  T_1286;
  wire [7:0] T_1290;
  wire [7:0] T_1294;
  wire [7:0] T_1298;
  wire [7:0] T_1302;
  wire [7:0] T_1306;
  wire [7:0] T_1310;
  wire [7:0] T_1314;
  wire [7:0] T_1318;
  wire [15:0] T_1319;
  wire [15:0] T_1320;
  wire [31:0] T_1321;
  wire [15:0] T_1322;
  wire [15:0] T_1323;
  wire [31:0] T_1324;
  wire [63:0] T_1325;
  wire [63:0] T_1326;
  wire [63:0] T_1403;
  wire [63:0] T_1404;
  wire [63:0] masked_wdata;
  wire  T_1406;
  wire [35:0] T_1409;
  wire  GEN_1;
  wire [36:0] T_1410;
  wire [7:0] T_1412;
  wire [36:0] T_1413;
  wire  T_1414;
  wire  T_1415;
  wire  GEN_2;
  wire  GEN_101;
  wire  GEN_102;
  wire  GEN_103;
  wire  GEN_104;
  wire  GEN_105;
  wire  GEN_106;
  wire  GEN_107;
  wire  GEN_108;
  wire  GEN_109;
  wire  GEN_110;
  wire  GEN_111;
  wire  GEN_112;
  wire  GEN_113;
  wire  GEN_114;
  wire  GEN_115;
  wire  GEN_116;
  wire  GEN_117;
  wire  GEN_118;
  wire  GEN_119;
  wire  GEN_120;
  wire  GEN_121;
  wire  GEN_122;
  wire  GEN_123;
  wire  GEN_124;
  wire  GEN_125;
  wire  GEN_126;
  wire  GEN_127;
  wire  GEN_128;
  wire  GEN_129;
  wire  GEN_130;
  wire  GEN_131;
  wire  GEN_134;
  wire  GEN_135;
  wire  GEN_136;
  wire  GEN_137;
  wire  GEN_138;
  wire  GEN_139;
  wire  GEN_140;
  wire  GEN_141;
  wire  GEN_142;
  wire  GEN_143;
  wire  GEN_144;
  wire  GEN_145;
  wire  GEN_146;
  wire  GEN_147;
  wire  GEN_148;
  wire  GEN_149;
  wire  GEN_150;
  wire  GEN_151;
  wire  GEN_152;
  wire  GEN_153;
  wire  GEN_154;
  wire  GEN_155;
  wire  GEN_156;
  wire  GEN_157;
  wire  GEN_158;
  wire  GEN_159;
  wire  GEN_160;
  wire  GEN_161;
  wire  GEN_162;
  wire  GEN_163;
  wire  GEN_164;
  wire [31:0] T_1447;
  wire [4:0] T_1448;
  wire  GEN_3;
  wire  GEN_717;
  wire  GEN_718;
  wire  GEN_165;
  wire  GEN_720;
  wire  GEN_166;
  wire  GEN_722;
  wire  GEN_167;
  wire  GEN_724;
  wire  GEN_168;
  wire  GEN_726;
  wire  GEN_169;
  wire  GEN_728;
  wire  GEN_170;
  wire  GEN_730;
  wire  GEN_171;
  wire  GEN_732;
  wire  GEN_172;
  wire  GEN_734;
  wire  GEN_173;
  wire  GEN_736;
  wire  GEN_174;
  wire  GEN_738;
  wire  GEN_175;
  wire  GEN_740;
  wire  GEN_176;
  wire  GEN_742;
  wire  GEN_177;
  wire  GEN_744;
  wire  GEN_178;
  wire  GEN_746;
  wire  GEN_179;
  wire  GEN_748;
  wire  GEN_180;
  wire  GEN_750;
  wire  GEN_181;
  wire  GEN_752;
  wire  GEN_182;
  wire  GEN_754;
  wire  GEN_183;
  wire  GEN_756;
  wire  GEN_184;
  wire  GEN_758;
  wire  GEN_185;
  wire  GEN_760;
  wire  GEN_186;
  wire  GEN_762;
  wire  GEN_187;
  wire  GEN_764;
  wire  GEN_188;
  wire  GEN_766;
  wire  GEN_189;
  wire  GEN_768;
  wire  GEN_190;
  wire  GEN_770;
  wire  GEN_191;
  wire  GEN_772;
  wire  GEN_192;
  wire  GEN_774;
  wire  GEN_193;
  wire  GEN_776;
  wire  GEN_194;
  wire  GEN_778;
  wire  GEN_195;
  wire [5:0] T_1450;
  wire [4:0] T_1451;
  wire  GEN_4;
  wire  GEN_196;
  wire  GEN_197;
  wire  GEN_198;
  wire  GEN_199;
  wire  GEN_200;
  wire  GEN_201;
  wire  GEN_202;
  wire  GEN_203;
  wire  GEN_204;
  wire  GEN_205;
  wire  GEN_206;
  wire  GEN_207;
  wire  GEN_208;
  wire  GEN_209;
  wire  GEN_210;
  wire  GEN_211;
  wire  GEN_212;
  wire  GEN_213;
  wire  GEN_214;
  wire  GEN_215;
  wire  GEN_216;
  wire  GEN_217;
  wire  GEN_218;
  wire  GEN_219;
  wire  GEN_220;
  wire  GEN_221;
  wire  GEN_222;
  wire  GEN_223;
  wire  GEN_224;
  wire  GEN_225;
  wire  GEN_226;
  wire  GEN_228;
  wire  GEN_229;
  wire  GEN_230;
  wire  GEN_231;
  wire  GEN_232;
  wire  GEN_233;
  wire  GEN_234;
  wire  GEN_235;
  wire  GEN_236;
  wire  GEN_237;
  wire  GEN_238;
  wire  GEN_239;
  wire  GEN_240;
  wire  GEN_241;
  wire  GEN_242;
  wire  GEN_243;
  wire  GEN_244;
  wire  GEN_245;
  wire  GEN_246;
  wire  GEN_247;
  wire  GEN_248;
  wire  GEN_249;
  wire  GEN_250;
  wire  GEN_251;
  wire  GEN_252;
  wire  GEN_253;
  wire  GEN_254;
  wire  GEN_255;
  wire  GEN_256;
  wire  GEN_257;
  wire  GEN_258;
  wire  GEN_261;
  wire  GEN_262;
  wire  GEN_263;
  wire  GEN_264;
  wire  GEN_265;
  wire  GEN_266;
  wire  GEN_267;
  wire  GEN_268;
  wire  GEN_269;
  wire  GEN_270;
  wire  GEN_271;
  wire  GEN_272;
  wire  GEN_273;
  wire  GEN_274;
  wire  GEN_275;
  wire  GEN_276;
  wire  GEN_277;
  wire  GEN_278;
  wire  GEN_279;
  wire  GEN_280;
  wire  GEN_281;
  wire  GEN_282;
  wire  GEN_283;
  wire  GEN_284;
  wire  GEN_285;
  wire  GEN_286;
  wire  GEN_287;
  wire  GEN_288;
  wire  GEN_289;
  wire  GEN_290;
  wire  GEN_291;
  wire  GEN_294;
  wire  GEN_295;
  wire  GEN_296;
  wire  GEN_297;
  wire  GEN_298;
  wire  GEN_299;
  wire  GEN_300;
  wire  GEN_301;
  wire  GEN_302;
  wire  GEN_303;
  wire  GEN_304;
  wire  GEN_305;
  wire  GEN_306;
  wire  GEN_307;
  wire  GEN_308;
  wire  GEN_309;
  wire  GEN_310;
  wire  GEN_311;
  wire  GEN_312;
  wire  GEN_313;
  wire  GEN_314;
  wire  GEN_315;
  wire  GEN_316;
  wire  GEN_317;
  wire  GEN_318;
  wire  GEN_319;
  wire  GEN_320;
  wire  GEN_321;
  wire  GEN_322;
  wire  GEN_323;
  wire  GEN_324;
  wire [63:0] GEN_326;
  wire  GEN_329;
  wire  GEN_330;
  wire  GEN_331;
  wire  GEN_332;
  wire  GEN_333;
  wire  GEN_334;
  wire  GEN_335;
  wire  GEN_336;
  wire  GEN_337;
  wire  GEN_338;
  wire  GEN_339;
  wire  GEN_340;
  wire  GEN_341;
  wire  GEN_342;
  wire  GEN_343;
  wire  GEN_344;
  wire  GEN_345;
  wire  GEN_346;
  wire  GEN_347;
  wire  GEN_348;
  wire  GEN_349;
  wire  GEN_350;
  wire  GEN_351;
  wire  GEN_352;
  wire  GEN_353;
  wire  GEN_354;
  wire  GEN_355;
  wire  GEN_356;
  wire  GEN_357;
  wire  GEN_358;
  wire  GEN_359;
  wire  GEN_362;
  wire  GEN_363;
  wire  GEN_364;
  wire  GEN_365;
  wire  GEN_366;
  wire  GEN_367;
  wire  GEN_368;
  wire  GEN_369;
  wire  GEN_370;
  wire  GEN_371;
  wire  GEN_372;
  wire  GEN_373;
  wire  GEN_374;
  wire  GEN_375;
  wire  GEN_376;
  wire  GEN_377;
  wire  GEN_378;
  wire  GEN_379;
  wire  GEN_380;
  wire  GEN_381;
  wire  GEN_382;
  wire  GEN_383;
  wire  GEN_384;
  wire  GEN_385;
  wire  GEN_386;
  wire  GEN_387;
  wire  GEN_388;
  wire  GEN_389;
  wire  GEN_390;
  wire  GEN_391;
  wire  GEN_392;
  wire  T_1459;
  wire  T_1461;
  wire  T_1462;
  wire  GEN_5;
  wire  GEN_6;
  wire [1:0] T_1467;
  wire  GEN_7;
  wire  GEN_8;
  wire [1:0] T_1468;
  wire [3:0] T_1469;
  wire  GEN_9;
  wire  GEN_10;
  wire [1:0] T_1470;
  wire  GEN_11;
  wire  GEN_12;
  wire [1:0] T_1471;
  wire [3:0] T_1472;
  wire [7:0] T_1473;
  wire  GEN_13;
  wire  GEN_14;
  wire [1:0] T_1474;
  wire  GEN_15;
  wire  GEN_16;
  wire [1:0] T_1475;
  wire [3:0] T_1476;
  wire  GEN_17;
  wire  GEN_18;
  wire [1:0] T_1477;
  wire  GEN_19;
  wire  GEN_20;
  wire [1:0] T_1478;
  wire [3:0] T_1479;
  wire [7:0] T_1480;
  wire [15:0] T_1481;
  wire  GEN_21;
  wire  GEN_22;
  wire [1:0] T_1482;
  wire  GEN_23;
  wire  GEN_24;
  wire [1:0] T_1483;
  wire [3:0] T_1484;
  wire  GEN_25;
  wire  GEN_26;
  wire [1:0] T_1485;
  wire  GEN_27;
  wire  GEN_28;
  wire [1:0] T_1486;
  wire [3:0] T_1487;
  wire [7:0] T_1488;
  wire  GEN_29;
  wire  GEN_30;
  wire [1:0] T_1489;
  wire  GEN_31;
  wire  GEN_32;
  wire [1:0] T_1490;
  wire [3:0] T_1491;
  wire  GEN_33;
  wire  GEN_34;
  wire [1:0] T_1492;
  wire  GEN_35;
  wire  GEN_36;
  wire [1:0] T_1493;
  wire [3:0] T_1494;
  wire [7:0] T_1495;
  wire [15:0] T_1496;
  wire [31:0] T_1497;
  wire  T_1501;
  wire  GEN_37;
  wire  T_1505;
  wire  GEN_38;
  wire  GEN_398;
  wire  T_1509;
  wire  GEN_39;
  wire  GEN_401;
  wire  T_1513;
  wire  GEN_40;
  wire  GEN_404;
  wire  T_1517;
  wire  GEN_41;
  wire  GEN_407;
  wire  T_1521;
  wire  GEN_42;
  wire  GEN_410;
  wire  T_1525;
  wire  GEN_43;
  wire  GEN_413;
  wire  T_1529;
  wire  GEN_44;
  wire  GEN_416;
  wire  T_1533;
  wire  GEN_45;
  wire  GEN_419;
  wire  T_1537;
  wire  GEN_46;
  wire  GEN_422;
  wire  T_1541;
  wire  GEN_47;
  wire  GEN_425;
  wire  T_1545;
  wire  GEN_48;
  wire  GEN_428;
  wire  T_1549;
  wire  GEN_49;
  wire  GEN_431;
  wire  T_1553;
  wire  GEN_50;
  wire  GEN_434;
  wire  T_1557;
  wire  GEN_51;
  wire  GEN_437;
  wire  T_1561;
  wire  GEN_52;
  wire  GEN_440;
  wire  T_1565;
  wire  GEN_53;
  wire  GEN_443;
  wire  T_1569;
  wire  GEN_54;
  wire  GEN_446;
  wire  T_1573;
  wire  GEN_55;
  wire  GEN_449;
  wire  T_1577;
  wire  GEN_56;
  wire  GEN_452;
  wire  T_1581;
  wire  GEN_57;
  wire  GEN_455;
  wire  T_1585;
  wire  GEN_58;
  wire  GEN_458;
  wire  T_1589;
  wire  GEN_59;
  wire  GEN_461;
  wire  T_1593;
  wire  GEN_60;
  wire  GEN_464;
  wire  T_1597;
  wire  GEN_61;
  wire  GEN_467;
  wire  T_1601;
  wire  GEN_62;
  wire  GEN_470;
  wire  T_1605;
  wire  GEN_63;
  wire  GEN_473;
  wire  T_1609;
  wire  GEN_64;
  wire  GEN_476;
  wire  T_1613;
  wire  GEN_65;
  wire  GEN_479;
  wire  T_1617;
  wire  GEN_66;
  wire  GEN_482;
  wire  T_1621;
  wire  GEN_67;
  wire  GEN_485;
  wire  T_1625;
  wire  GEN_68;
  wire  GEN_488;
  wire [63:0] GEN_521;
  wire [63:0] GEN_619;
  wire  GEN_623;
  wire  GEN_625;
  wire  GEN_627;
  wire  GEN_629;
  wire  GEN_631;
  wire  GEN_633;
  wire  GEN_635;
  wire  GEN_637;
  wire  GEN_639;
  wire  GEN_641;
  wire  GEN_643;
  wire  GEN_645;
  wire  GEN_647;
  wire  GEN_649;
  wire  GEN_651;
  wire  GEN_653;
  wire  GEN_655;
  wire  GEN_657;
  wire  GEN_659;
  wire  GEN_661;
  wire  GEN_663;
  wire  GEN_665;
  wire  GEN_667;
  wire  GEN_669;
  wire  GEN_671;
  wire  GEN_673;
  wire  GEN_675;
  wire  GEN_677;
  wire  GEN_679;
  wire  GEN_681;
  wire  GEN_683;
  wire  T_1627;
  wire  T_1631;
  wire  T_1632;
  wire  T_1633;
  wire [1:0] T_1634;
  wire [1:0] T_1635;
  wire [1:0] T_1636;
  wire [3:0] T_1637;
  wire [1:0] T_1638;
  wire [1:0] T_1639;
  wire [3:0] T_1640;
  wire [7:0] T_1641;
  wire [1:0] T_1642;
  wire [1:0] T_1643;
  wire [3:0] T_1644;
  wire [1:0] T_1645;
  wire [1:0] T_1646;
  wire [3:0] T_1647;
  wire [7:0] T_1648;
  wire [15:0] T_1649;
  wire [1:0] T_1650;
  wire [1:0] T_1651;
  wire [3:0] T_1652;
  wire [1:0] T_1653;
  wire [1:0] T_1654;
  wire [3:0] T_1655;
  wire [7:0] T_1656;
  wire [1:0] T_1657;
  wire [1:0] T_1658;
  wire [3:0] T_1659;
  wire [1:0] T_1660;
  wire [1:0] T_1661;
  wire [3:0] T_1662;
  wire [7:0] T_1663;
  wire [15:0] T_1664;
  wire [31:0] T_1665;
  wire [6:0] GEN_779;
  wire [8:0] T_1667;
  wire [31:0] T_1668;
  wire [63:0] GEN_684;
  wire  T_1675;
  wire  T_1676;
  wire [3:0] T_1677;
  wire  T_1679;
  wire [31:0] T_1681;
  wire [31:0] T_1683;
  wire [63:0] T_1684;
  wire [63:0] GEN_685;
  wire  T_1686;
  wire [31:0] T_1688;
  wire [31:0] T_1690;
  wire [63:0] T_1691;
  wire [63:0] GEN_686;
  wire  T_1693;
  wire [31:0] T_1695;
  wire [31:0] T_1697;
  wire [63:0] T_1698;
  wire [63:0] GEN_687;
  wire  T_1700;
  wire [31:0] T_1702;
  wire [31:0] T_1704;
  wire [63:0] T_1705;
  wire [63:0] GEN_688;
  wire  T_1707;
  wire [31:0] T_1709;
  wire [31:0] T_1711;
  wire [63:0] T_1712;
  wire [63:0] GEN_689;
  wire  T_1714;
  wire [31:0] T_1716;
  wire [31:0] T_1718;
  wire [63:0] T_1719;
  wire [63:0] GEN_690;
  wire  T_1721;
  wire [31:0] T_1723;
  wire [31:0] T_1725;
  wire [63:0] T_1726;
  wire [63:0] GEN_691;
  wire  T_1728;
  wire [31:0] T_1730;
  wire [31:0] T_1732;
  wire [63:0] T_1733;
  wire [63:0] GEN_692;
  wire  T_1735;
  wire [31:0] T_1737;
  wire [31:0] T_1739;
  wire [63:0] T_1740;
  wire [63:0] GEN_693;
  wire  T_1742;
  wire [31:0] T_1744;
  wire [31:0] T_1746;
  wire [63:0] T_1747;
  wire [63:0] GEN_694;
  wire  T_1749;
  wire [31:0] T_1751;
  wire [31:0] T_1753;
  wire [63:0] T_1754;
  wire [63:0] GEN_695;
  wire  T_1756;
  wire [31:0] T_1758;
  wire [31:0] T_1760;
  wire [63:0] T_1761;
  wire [63:0] GEN_696;
  wire  T_1763;
  wire [31:0] T_1765;
  wire [31:0] T_1767;
  wire [63:0] T_1768;
  wire [63:0] GEN_697;
  wire  T_1770;
  wire [31:0] T_1772;
  wire [31:0] T_1774;
  wire [63:0] T_1775;
  wire [63:0] GEN_698;
  wire  T_1777;
  wire [31:0] T_1779;
  wire [31:0] T_1781;
  wire [63:0] T_1782;
  wire [63:0] GEN_699;
  wire  T_1784;
  wire [31:0] T_1786;
  wire [31:0] T_1788;
  wire [63:0] T_1789;
  wire [63:0] GEN_700;
  wire [63:0] GEN_701;
  wire  T_1809;
  wire [2:0] T_1810;
  wire  T_1811;
  wire [2:0] T_1812;
  wire  T_1813;
  wire [2:0] T_1814;
  wire  T_1815;
  wire [2:0] T_1816;
  wire  T_1817;
  wire [2:0] T_1818;
  wire  T_1819;
  wire [2:0] T_1820;
  wire  T_1821;
  wire [2:0] T_1822;
  wire [2:0] T_1847_addr_beat;
  wire [1:0] T_1847_client_xact_id;
  wire  T_1847_manager_xact_id;
  wire  T_1847_is_builtin_type;
  wire [3:0] T_1847_g_type;
  wire [63:0] T_1847_data;
  Queue_8 acq (
    .clk(acq_clk),
    .reset(acq_reset),
    .io_enq_ready(acq_io_enq_ready),
    .io_enq_valid(acq_io_enq_valid),
    .io_enq_bits_addr_block(acq_io_enq_bits_addr_block),
    .io_enq_bits_client_xact_id(acq_io_enq_bits_client_xact_id),
    .io_enq_bits_addr_beat(acq_io_enq_bits_addr_beat),
    .io_enq_bits_is_builtin_type(acq_io_enq_bits_is_builtin_type),
    .io_enq_bits_a_type(acq_io_enq_bits_a_type),
    .io_enq_bits_union(acq_io_enq_bits_union),
    .io_enq_bits_data(acq_io_enq_bits_data),
    .io_deq_ready(acq_io_deq_ready),
    .io_deq_valid(acq_io_deq_valid),
    .io_deq_bits_addr_block(acq_io_deq_bits_addr_block),
    .io_deq_bits_client_xact_id(acq_io_deq_bits_client_xact_id),
    .io_deq_bits_addr_beat(acq_io_deq_bits_addr_beat),
    .io_deq_bits_is_builtin_type(acq_io_deq_bits_is_builtin_type),
    .io_deq_bits_a_type(acq_io_deq_bits_a_type),
    .io_deq_bits_union(acq_io_deq_bits_union),
    .io_deq_bits_data(acq_io_deq_bits_data),
    .io_count(acq_io_count)
  );
  assign io_devices_0_ready = T_770;
  assign io_devices_0_complete = GEN_362;
  assign io_devices_1_ready = T_774;
  assign io_devices_1_complete = GEN_363;
  assign io_devices_2_ready = T_778;
  assign io_devices_2_complete = GEN_364;
  assign io_devices_3_ready = T_782;
  assign io_devices_3_complete = GEN_365;
  assign io_devices_4_ready = T_786;
  assign io_devices_4_complete = GEN_366;
  assign io_devices_5_ready = T_790;
  assign io_devices_5_complete = GEN_367;
  assign io_devices_6_ready = T_794;
  assign io_devices_6_complete = GEN_368;
  assign io_devices_7_ready = T_798;
  assign io_devices_7_complete = GEN_369;
  assign io_devices_8_ready = T_802;
  assign io_devices_8_complete = GEN_370;
  assign io_devices_9_ready = T_806;
  assign io_devices_9_complete = GEN_371;
  assign io_devices_10_ready = T_810;
  assign io_devices_10_complete = GEN_372;
  assign io_devices_11_ready = T_814;
  assign io_devices_11_complete = GEN_373;
  assign io_devices_12_ready = T_818;
  assign io_devices_12_complete = GEN_374;
  assign io_devices_13_ready = T_822;
  assign io_devices_13_complete = GEN_375;
  assign io_devices_14_ready = T_826;
  assign io_devices_14_complete = GEN_376;
  assign io_devices_15_ready = T_830;
  assign io_devices_15_complete = GEN_377;
  assign io_devices_16_ready = T_834;
  assign io_devices_16_complete = GEN_378;
  assign io_devices_17_ready = T_838;
  assign io_devices_17_complete = GEN_379;
  assign io_devices_18_ready = T_842;
  assign io_devices_18_complete = GEN_380;
  assign io_devices_19_ready = T_846;
  assign io_devices_19_complete = GEN_381;
  assign io_devices_20_ready = T_850;
  assign io_devices_20_complete = GEN_382;
  assign io_devices_21_ready = T_854;
  assign io_devices_21_complete = GEN_383;
  assign io_devices_22_ready = T_858;
  assign io_devices_22_complete = GEN_384;
  assign io_devices_23_ready = T_862;
  assign io_devices_23_complete = GEN_385;
  assign io_devices_24_ready = T_866;
  assign io_devices_24_complete = GEN_386;
  assign io_devices_25_ready = T_870;
  assign io_devices_25_complete = GEN_387;
  assign io_devices_26_ready = T_874;
  assign io_devices_26_complete = GEN_388;
  assign io_devices_27_ready = T_878;
  assign io_devices_27_complete = GEN_389;
  assign io_devices_28_ready = T_882;
  assign io_devices_28_complete = GEN_390;
  assign io_devices_29_ready = T_886;
  assign io_devices_29_complete = GEN_391;
  assign io_devices_30_ready = T_890;
  assign io_devices_30_complete = GEN_392;
  assign io_harts_0 = T_1186;
  assign io_tl_acquire_ready = acq_io_enq_ready;
  assign io_tl_grant_valid = acq_io_deq_valid;
  assign io_tl_grant_bits_addr_beat = T_1847_addr_beat;
  assign io_tl_grant_bits_client_xact_id = T_1847_client_xact_id;
  assign io_tl_grant_bits_manager_xact_id = T_1847_manager_xact_id;
  assign io_tl_grant_bits_is_builtin_type = T_1847_is_builtin_type;
  assign io_tl_grant_bits_g_type = T_1847_g_type;
  assign io_tl_grant_bits_data = T_1847_data;
  assign T_680_0 = 1'h1;
  assign T_680_1 = 1'h1;
  assign T_680_2 = 1'h1;
  assign T_680_3 = 1'h1;
  assign T_680_4 = 1'h1;
  assign T_680_5 = 1'h1;
  assign T_680_6 = 1'h1;
  assign T_680_7 = 1'h1;
  assign T_680_8 = 1'h1;
  assign T_680_9 = 1'h1;
  assign T_680_10 = 1'h1;
  assign T_680_11 = 1'h1;
  assign T_680_12 = 1'h1;
  assign T_680_13 = 1'h1;
  assign T_680_14 = 1'h1;
  assign T_680_15 = 1'h1;
  assign T_680_16 = 1'h1;
  assign T_680_17 = 1'h1;
  assign T_680_18 = 1'h1;
  assign T_680_19 = 1'h1;
  assign T_680_20 = 1'h1;
  assign T_680_21 = 1'h1;
  assign T_680_22 = 1'h1;
  assign T_680_23 = 1'h1;
  assign T_680_24 = 1'h1;
  assign T_680_25 = 1'h1;
  assign T_680_26 = 1'h1;
  assign T_680_27 = 1'h1;
  assign T_680_28 = 1'h1;
  assign T_680_29 = 1'h1;
  assign T_680_30 = 1'h1;
  assign T_680_31 = 1'h1;
  assign priority_0 = 1'h0;
  assign priority_1 = T_680_1;
  assign priority_2 = T_680_2;
  assign priority_3 = T_680_3;
  assign priority_4 = T_680_4;
  assign priority_5 = T_680_5;
  assign priority_6 = T_680_6;
  assign priority_7 = T_680_7;
  assign priority_8 = T_680_8;
  assign priority_9 = T_680_9;
  assign priority_10 = T_680_10;
  assign priority_11 = T_680_11;
  assign priority_12 = T_680_12;
  assign priority_13 = T_680_13;
  assign priority_14 = T_680_14;
  assign priority_15 = T_680_15;
  assign priority_16 = T_680_16;
  assign priority_17 = T_680_17;
  assign priority_18 = T_680_18;
  assign priority_19 = T_680_19;
  assign priority_20 = T_680_20;
  assign priority_21 = T_680_21;
  assign priority_22 = T_680_22;
  assign priority_23 = T_680_23;
  assign priority_24 = T_680_24;
  assign priority_25 = T_680_25;
  assign priority_26 = T_680_26;
  assign priority_27 = T_680_27;
  assign priority_28 = T_680_28;
  assign priority_29 = T_680_29;
  assign priority_30 = T_680_30;
  assign priority_31 = T_680_31;
  assign T_691_0 = 1'h0;
  assign threshold_0 = T_691_0;
  assign T_733_0 = 1'h0;
  assign T_733_1 = 1'h0;
  assign T_733_2 = 1'h0;
  assign T_733_3 = 1'h0;
  assign T_733_4 = 1'h0;
  assign T_733_5 = 1'h0;
  assign T_733_6 = 1'h0;
  assign T_733_7 = 1'h0;
  assign T_733_8 = 1'h0;
  assign T_733_9 = 1'h0;
  assign T_733_10 = 1'h0;
  assign T_733_11 = 1'h0;
  assign T_733_12 = 1'h0;
  assign T_733_13 = 1'h0;
  assign T_733_14 = 1'h0;
  assign T_733_15 = 1'h0;
  assign T_733_16 = 1'h0;
  assign T_733_17 = 1'h0;
  assign T_733_18 = 1'h0;
  assign T_733_19 = 1'h0;
  assign T_733_20 = 1'h0;
  assign T_733_21 = 1'h0;
  assign T_733_22 = 1'h0;
  assign T_733_23 = 1'h0;
  assign T_733_24 = 1'h0;
  assign T_733_25 = 1'h0;
  assign T_733_26 = 1'h0;
  assign T_733_27 = 1'h0;
  assign T_733_28 = 1'h0;
  assign T_733_29 = 1'h0;
  assign T_733_30 = 1'h0;
  assign T_733_31 = 1'h0;
  assign T_770 = pending_1 == 1'h0;
  assign GEN_69 = io_devices_0_valid ? 1'h1 : pending_1;
  assign T_774 = pending_2 == 1'h0;
  assign GEN_70 = io_devices_1_valid ? 1'h1 : pending_2;
  assign T_778 = pending_3 == 1'h0;
  assign GEN_71 = io_devices_2_valid ? 1'h1 : pending_3;
  assign T_782 = pending_4 == 1'h0;
  assign GEN_72 = io_devices_3_valid ? 1'h1 : pending_4;
  assign T_786 = pending_5 == 1'h0;
  assign GEN_73 = io_devices_4_valid ? 1'h1 : pending_5;
  assign T_790 = pending_6 == 1'h0;
  assign GEN_74 = io_devices_5_valid ? 1'h1 : pending_6;
  assign T_794 = pending_7 == 1'h0;
  assign GEN_75 = io_devices_6_valid ? 1'h1 : pending_7;
  assign T_798 = pending_8 == 1'h0;
  assign GEN_76 = io_devices_7_valid ? 1'h1 : pending_8;
  assign T_802 = pending_9 == 1'h0;
  assign GEN_77 = io_devices_8_valid ? 1'h1 : pending_9;
  assign T_806 = pending_10 == 1'h0;
  assign GEN_78 = io_devices_9_valid ? 1'h1 : pending_10;
  assign T_810 = pending_11 == 1'h0;
  assign GEN_79 = io_devices_10_valid ? 1'h1 : pending_11;
  assign T_814 = pending_12 == 1'h0;
  assign GEN_80 = io_devices_11_valid ? 1'h1 : pending_12;
  assign T_818 = pending_13 == 1'h0;
  assign GEN_81 = io_devices_12_valid ? 1'h1 : pending_13;
  assign T_822 = pending_14 == 1'h0;
  assign GEN_82 = io_devices_13_valid ? 1'h1 : pending_14;
  assign T_826 = pending_15 == 1'h0;
  assign GEN_83 = io_devices_14_valid ? 1'h1 : pending_15;
  assign T_830 = pending_16 == 1'h0;
  assign GEN_84 = io_devices_15_valid ? 1'h1 : pending_16;
  assign T_834 = pending_17 == 1'h0;
  assign GEN_85 = io_devices_16_valid ? 1'h1 : pending_17;
  assign T_838 = pending_18 == 1'h0;
  assign GEN_86 = io_devices_17_valid ? 1'h1 : pending_18;
  assign T_842 = pending_19 == 1'h0;
  assign GEN_87 = io_devices_18_valid ? 1'h1 : pending_19;
  assign T_846 = pending_20 == 1'h0;
  assign GEN_88 = io_devices_19_valid ? 1'h1 : pending_20;
  assign T_850 = pending_21 == 1'h0;
  assign GEN_89 = io_devices_20_valid ? 1'h1 : pending_21;
  assign T_854 = pending_22 == 1'h0;
  assign GEN_90 = io_devices_21_valid ? 1'h1 : pending_22;
  assign T_858 = pending_23 == 1'h0;
  assign GEN_91 = io_devices_22_valid ? 1'h1 : pending_23;
  assign T_862 = pending_24 == 1'h0;
  assign GEN_92 = io_devices_23_valid ? 1'h1 : pending_24;
  assign T_866 = pending_25 == 1'h0;
  assign GEN_93 = io_devices_24_valid ? 1'h1 : pending_25;
  assign T_870 = pending_26 == 1'h0;
  assign GEN_94 = io_devices_25_valid ? 1'h1 : pending_26;
  assign T_874 = pending_27 == 1'h0;
  assign GEN_95 = io_devices_26_valid ? 1'h1 : pending_27;
  assign T_878 = pending_28 == 1'h0;
  assign GEN_96 = io_devices_27_valid ? 1'h1 : pending_28;
  assign T_882 = pending_29 == 1'h0;
  assign GEN_97 = io_devices_28_valid ? 1'h1 : pending_29;
  assign T_886 = pending_30 == 1'h0;
  assign GEN_98 = io_devices_29_valid ? 1'h1 : pending_30;
  assign T_890 = pending_31 == 1'h0;
  assign GEN_99 = io_devices_30_valid ? 1'h1 : pending_31;
  assign maxDevs_0 = T_1182;
  assign T_900 = pending_1 & enables_0_1;
  assign T_901 = {T_900,priority_1};
  assign T_902 = pending_2 & enables_0_2;
  assign T_903 = {T_902,priority_2};
  assign T_904 = pending_3 & enables_0_3;
  assign T_905 = {T_904,priority_3};
  assign T_906 = pending_4 & enables_0_4;
  assign T_907 = {T_906,priority_4};
  assign T_908 = pending_5 & enables_0_5;
  assign T_909 = {T_908,priority_5};
  assign T_910 = pending_6 & enables_0_6;
  assign T_911 = {T_910,priority_6};
  assign T_912 = pending_7 & enables_0_7;
  assign T_913 = {T_912,priority_7};
  assign T_914 = pending_8 & enables_0_8;
  assign T_915 = {T_914,priority_8};
  assign T_916 = pending_9 & enables_0_9;
  assign T_917 = {T_916,priority_9};
  assign T_918 = pending_10 & enables_0_10;
  assign T_919 = {T_918,priority_10};
  assign T_920 = pending_11 & enables_0_11;
  assign T_921 = {T_920,priority_11};
  assign T_922 = pending_12 & enables_0_12;
  assign T_923 = {T_922,priority_12};
  assign T_924 = pending_13 & enables_0_13;
  assign T_925 = {T_924,priority_13};
  assign T_926 = pending_14 & enables_0_14;
  assign T_927 = {T_926,priority_14};
  assign T_928 = pending_15 & enables_0_15;
  assign T_929 = {T_928,priority_15};
  assign T_930 = pending_16 & enables_0_16;
  assign T_931 = {T_930,priority_16};
  assign T_932 = pending_17 & enables_0_17;
  assign T_933 = {T_932,priority_17};
  assign T_934 = pending_18 & enables_0_18;
  assign T_935 = {T_934,priority_18};
  assign T_936 = pending_19 & enables_0_19;
  assign T_937 = {T_936,priority_19};
  assign T_938 = pending_20 & enables_0_20;
  assign T_939 = {T_938,priority_20};
  assign T_940 = pending_21 & enables_0_21;
  assign T_941 = {T_940,priority_21};
  assign T_942 = pending_22 & enables_0_22;
  assign T_943 = {T_942,priority_22};
  assign T_944 = pending_23 & enables_0_23;
  assign T_945 = {T_944,priority_23};
  assign T_946 = pending_24 & enables_0_24;
  assign T_947 = {T_946,priority_24};
  assign T_948 = pending_25 & enables_0_25;
  assign T_949 = {T_948,priority_25};
  assign T_950 = pending_26 & enables_0_26;
  assign T_951 = {T_950,priority_26};
  assign T_952 = pending_27 & enables_0_27;
  assign T_953 = {T_952,priority_27};
  assign T_954 = pending_28 & enables_0_28;
  assign T_955 = {T_954,priority_28};
  assign T_956 = pending_29 & enables_0_29;
  assign T_957 = {T_956,priority_29};
  assign T_958 = pending_30 & enables_0_30;
  assign T_959 = {T_958,priority_30};
  assign T_960 = pending_31 & enables_0_31;
  assign T_961 = {T_960,priority_31};
  assign T_966 = 2'h2 >= T_901;
  assign T_967 = T_966 ? 2'h2 : T_901;
  assign T_969 = 1'h1 + 1'h0;
  assign T_970 = T_969[0:0];
  assign T_971 = T_966 ? 1'h0 : T_970;
  assign T_974 = T_903 >= T_905;
  assign T_975 = T_974 ? T_903 : T_905;
  assign T_979 = T_974 ? 1'h0 : T_970;
  assign T_980 = T_967 >= T_975;
  assign T_981 = T_980 ? T_967 : T_975;
  assign GEN_702 = {{1'd0}, T_979};
  assign T_983 = 2'h2 + GEN_702;
  assign T_984 = T_983[1:0];
  assign T_985 = T_980 ? {{1'd0}, T_971} : T_984;
  assign T_988 = T_907 >= T_909;
  assign T_989 = T_988 ? T_907 : T_909;
  assign T_993 = T_988 ? 1'h0 : T_970;
  assign T_996 = T_911 >= T_913;
  assign T_997 = T_996 ? T_911 : T_913;
  assign T_1001 = T_996 ? 1'h0 : T_970;
  assign T_1002 = T_989 >= T_997;
  assign T_1003 = T_1002 ? T_989 : T_997;
  assign GEN_703 = {{1'd0}, T_1001};
  assign T_1005 = 2'h2 + GEN_703;
  assign T_1006 = T_1005[1:0];
  assign T_1007 = T_1002 ? {{1'd0}, T_993} : T_1006;
  assign T_1008 = T_981 >= T_1003;
  assign T_1009 = T_1008 ? T_981 : T_1003;
  assign GEN_704 = {{1'd0}, T_1007};
  assign T_1011 = 3'h4 + GEN_704;
  assign T_1012 = T_1011[2:0];
  assign T_1013 = T_1008 ? {{1'd0}, T_985} : T_1012;
  assign T_1016 = T_915 >= T_917;
  assign T_1017 = T_1016 ? T_915 : T_917;
  assign T_1021 = T_1016 ? 1'h0 : T_970;
  assign T_1024 = T_919 >= T_921;
  assign T_1025 = T_1024 ? T_919 : T_921;
  assign T_1029 = T_1024 ? 1'h0 : T_970;
  assign T_1030 = T_1017 >= T_1025;
  assign T_1031 = T_1030 ? T_1017 : T_1025;
  assign GEN_705 = {{1'd0}, T_1029};
  assign T_1033 = 2'h2 + GEN_705;
  assign T_1034 = T_1033[1:0];
  assign T_1035 = T_1030 ? {{1'd0}, T_1021} : T_1034;
  assign T_1038 = T_923 >= T_925;
  assign T_1039 = T_1038 ? T_923 : T_925;
  assign T_1043 = T_1038 ? 1'h0 : T_970;
  assign T_1046 = T_927 >= T_929;
  assign T_1047 = T_1046 ? T_927 : T_929;
  assign T_1051 = T_1046 ? 1'h0 : T_970;
  assign T_1052 = T_1039 >= T_1047;
  assign T_1053 = T_1052 ? T_1039 : T_1047;
  assign GEN_706 = {{1'd0}, T_1051};
  assign T_1055 = 2'h2 + GEN_706;
  assign T_1056 = T_1055[1:0];
  assign T_1057 = T_1052 ? {{1'd0}, T_1043} : T_1056;
  assign T_1058 = T_1031 >= T_1053;
  assign T_1059 = T_1058 ? T_1031 : T_1053;
  assign GEN_707 = {{1'd0}, T_1057};
  assign T_1061 = 3'h4 + GEN_707;
  assign T_1062 = T_1061[2:0];
  assign T_1063 = T_1058 ? {{1'd0}, T_1035} : T_1062;
  assign T_1064 = T_1009 >= T_1059;
  assign T_1065 = T_1064 ? T_1009 : T_1059;
  assign GEN_708 = {{1'd0}, T_1063};
  assign T_1067 = 4'h8 + GEN_708;
  assign T_1068 = T_1067[3:0];
  assign T_1069 = T_1064 ? {{1'd0}, T_1013} : T_1068;
  assign T_1072 = T_931 >= T_933;
  assign T_1073 = T_1072 ? T_931 : T_933;
  assign T_1077 = T_1072 ? 1'h0 : T_970;
  assign T_1080 = T_935 >= T_937;
  assign T_1081 = T_1080 ? T_935 : T_937;
  assign T_1085 = T_1080 ? 1'h0 : T_970;
  assign T_1086 = T_1073 >= T_1081;
  assign T_1087 = T_1086 ? T_1073 : T_1081;
  assign GEN_709 = {{1'd0}, T_1085};
  assign T_1089 = 2'h2 + GEN_709;
  assign T_1090 = T_1089[1:0];
  assign T_1091 = T_1086 ? {{1'd0}, T_1077} : T_1090;
  assign T_1094 = T_939 >= T_941;
  assign T_1095 = T_1094 ? T_939 : T_941;
  assign T_1099 = T_1094 ? 1'h0 : T_970;
  assign T_1102 = T_943 >= T_945;
  assign T_1103 = T_1102 ? T_943 : T_945;
  assign T_1107 = T_1102 ? 1'h0 : T_970;
  assign T_1108 = T_1095 >= T_1103;
  assign T_1109 = T_1108 ? T_1095 : T_1103;
  assign GEN_710 = {{1'd0}, T_1107};
  assign T_1111 = 2'h2 + GEN_710;
  assign T_1112 = T_1111[1:0];
  assign T_1113 = T_1108 ? {{1'd0}, T_1099} : T_1112;
  assign T_1114 = T_1087 >= T_1109;
  assign T_1115 = T_1114 ? T_1087 : T_1109;
  assign GEN_711 = {{1'd0}, T_1113};
  assign T_1117 = 3'h4 + GEN_711;
  assign T_1118 = T_1117[2:0];
  assign T_1119 = T_1114 ? {{1'd0}, T_1091} : T_1118;
  assign T_1122 = T_947 >= T_949;
  assign T_1123 = T_1122 ? T_947 : T_949;
  assign T_1127 = T_1122 ? 1'h0 : T_970;
  assign T_1130 = T_951 >= T_953;
  assign T_1131 = T_1130 ? T_951 : T_953;
  assign T_1135 = T_1130 ? 1'h0 : T_970;
  assign T_1136 = T_1123 >= T_1131;
  assign T_1137 = T_1136 ? T_1123 : T_1131;
  assign GEN_712 = {{1'd0}, T_1135};
  assign T_1139 = 2'h2 + GEN_712;
  assign T_1140 = T_1139[1:0];
  assign T_1141 = T_1136 ? {{1'd0}, T_1127} : T_1140;
  assign T_1144 = T_955 >= T_957;
  assign T_1145 = T_1144 ? T_955 : T_957;
  assign T_1149 = T_1144 ? 1'h0 : T_970;
  assign T_1152 = T_959 >= T_961;
  assign T_1153 = T_1152 ? T_959 : T_961;
  assign T_1157 = T_1152 ? 1'h0 : T_970;
  assign T_1158 = T_1145 >= T_1153;
  assign T_1159 = T_1158 ? T_1145 : T_1153;
  assign GEN_713 = {{1'd0}, T_1157};
  assign T_1161 = 2'h2 + GEN_713;
  assign T_1162 = T_1161[1:0];
  assign T_1163 = T_1158 ? {{1'd0}, T_1149} : T_1162;
  assign T_1164 = T_1137 >= T_1159;
  assign T_1165 = T_1164 ? T_1137 : T_1159;
  assign GEN_714 = {{1'd0}, T_1163};
  assign T_1167 = 3'h4 + GEN_714;
  assign T_1168 = T_1167[2:0];
  assign T_1169 = T_1164 ? {{1'd0}, T_1141} : T_1168;
  assign T_1170 = T_1115 >= T_1165;
  assign T_1171 = T_1170 ? T_1115 : T_1165;
  assign GEN_715 = {{1'd0}, T_1169};
  assign T_1173 = 4'h8 + GEN_715;
  assign T_1174 = T_1173[3:0];
  assign T_1175 = T_1170 ? {{1'd0}, T_1119} : T_1174;
  assign T_1176 = T_1065 >= T_1171;
  assign T_1177 = T_1176 ? T_1065 : T_1171;
  assign GEN_716 = {{1'd0}, T_1175};
  assign T_1179 = 5'h10 + GEN_716;
  assign T_1180 = T_1179[4:0];
  assign T_1181 = T_1176 ? {{1'd0}, T_1069} : T_1180;
  assign T_1185 = {1'h1,threshold_0};
  assign T_1186 = T_1183 > T_1185;
  assign acq_clk = clk;
  assign acq_reset = reset;
  assign acq_io_enq_valid = io_tl_acquire_valid;
  assign acq_io_enq_bits_addr_block = io_tl_acquire_bits_addr_block;
  assign acq_io_enq_bits_client_xact_id = io_tl_acquire_bits_client_xact_id;
  assign acq_io_enq_bits_addr_beat = io_tl_acquire_bits_addr_beat;
  assign acq_io_enq_bits_is_builtin_type = io_tl_acquire_bits_is_builtin_type;
  assign acq_io_enq_bits_a_type = io_tl_acquire_bits_a_type;
  assign acq_io_enq_bits_union = io_tl_acquire_bits_union;
  assign acq_io_enq_bits_data = io_tl_acquire_bits_data;
  assign acq_io_deq_ready = io_tl_grant_ready;
  assign T_1210 = acq_io_deq_ready & acq_io_deq_valid;
  assign T_1212 = acq_io_deq_bits_a_type == 3'h0;
  assign T_1213 = acq_io_deq_bits_is_builtin_type & T_1212;
  assign read = T_1210 & T_1213;
  assign T_1216 = acq_io_deq_bits_a_type == 3'h2;
  assign T_1217 = acq_io_deq_bits_is_builtin_type & T_1216;
  assign write = T_1210 & T_1217;
  assign T_1220 = T_1210 == 1'h0;
  assign T_1221 = T_1220 | read;
  assign T_1222 = T_1221 | write;
  assign T_1223 = T_1222 | reset;
  assign T_1225 = T_1223 == 1'h0;
  assign T_1233_0 = 3'h0;
  assign T_1233_1 = 3'h4;
  assign T_1235 = acq_io_deq_bits_a_type == T_1233_0;
  assign T_1236 = acq_io_deq_bits_a_type == T_1233_1;
  assign T_1237 = T_1235 | T_1236;
  assign T_1238 = acq_io_deq_bits_is_builtin_type & T_1237;
  assign T_1239 = acq_io_deq_bits_union[11:9];
  assign T_1241 = T_1238 ? T_1239 : 3'h0;
  assign T_1242 = {acq_io_deq_bits_addr_block,acq_io_deq_bits_addr_beat};
  assign T_1243 = {T_1242,T_1241};
  assign addr = T_1243[25:0];
  assign hart = 1'h0;
  assign GEN_0 = maxDevs_0;
  assign T_1245 = GEN_0 + 5'h0;
  assign myMaxDev = T_1245[4:0];
  assign rdata = GEN_701;
  assign T_1251 = acq_io_deq_bits_a_type == 3'h4;
  assign T_1252 = acq_io_deq_bits_is_builtin_type & T_1251;
  assign T_1254 = T_1239[2];
  assign T_1256 = 2'h1 << T_1254;
  assign T_1257 = T_1256[0];
  assign T_1258 = T_1256[1];
  assign T_1262 = T_1257 ? 4'hf : 4'h0;
  assign T_1266 = T_1258 ? 4'hf : 4'h0;
  assign T_1267 = {T_1266,T_1262};
  assign T_1269 = acq_io_deq_bits_a_type == 3'h3;
  assign T_1270 = acq_io_deq_bits_is_builtin_type & T_1269;
  assign T_1274 = T_1270 | T_1217;
  assign T_1275 = acq_io_deq_bits_union[8:1];
  assign T_1277 = T_1274 ? T_1275 : 8'h0;
  assign T_1278 = T_1252 ? T_1267 : T_1277;
  assign T_1279 = T_1278[0];
  assign T_1280 = T_1278[1];
  assign T_1281 = T_1278[2];
  assign T_1282 = T_1278[3];
  assign T_1283 = T_1278[4];
  assign T_1284 = T_1278[5];
  assign T_1285 = T_1278[6];
  assign T_1286 = T_1278[7];
  assign T_1290 = T_1279 ? 8'hff : 8'h0;
  assign T_1294 = T_1280 ? 8'hff : 8'h0;
  assign T_1298 = T_1281 ? 8'hff : 8'h0;
  assign T_1302 = T_1282 ? 8'hff : 8'h0;
  assign T_1306 = T_1283 ? 8'hff : 8'h0;
  assign T_1310 = T_1284 ? 8'hff : 8'h0;
  assign T_1314 = T_1285 ? 8'hff : 8'h0;
  assign T_1318 = T_1286 ? 8'hff : 8'h0;
  assign T_1319 = {T_1294,T_1290};
  assign T_1320 = {T_1302,T_1298};
  assign T_1321 = {T_1320,T_1319};
  assign T_1322 = {T_1310,T_1306};
  assign T_1323 = {T_1318,T_1314};
  assign T_1324 = {T_1323,T_1322};
  assign T_1325 = {T_1324,T_1321};
  assign T_1326 = acq_io_deq_bits_data & T_1325;
  assign T_1403 = ~ T_1325;
  assign T_1404 = rdata & T_1403;
  assign masked_wdata = T_1326 | T_1404;
  assign T_1406 = addr >= 26'h200000;
  assign T_1409 = {myMaxDev,31'h0};
  assign GEN_1 = threshold_0;
  assign T_1410 = {T_1409,GEN_1};
  assign T_1412 = 7'h0 * 7'h40;
  assign T_1413 = T_1410 >> T_1412;
  assign T_1414 = addr[2];
  assign T_1415 = read & T_1414;
  assign GEN_2 = 1'h0;
  assign GEN_101 = 5'h1 == myMaxDev ? GEN_2 : GEN_69;
  assign GEN_102 = 5'h2 == myMaxDev ? GEN_2 : GEN_70;
  assign GEN_103 = 5'h3 == myMaxDev ? GEN_2 : GEN_71;
  assign GEN_104 = 5'h4 == myMaxDev ? GEN_2 : GEN_72;
  assign GEN_105 = 5'h5 == myMaxDev ? GEN_2 : GEN_73;
  assign GEN_106 = 5'h6 == myMaxDev ? GEN_2 : GEN_74;
  assign GEN_107 = 5'h7 == myMaxDev ? GEN_2 : GEN_75;
  assign GEN_108 = 5'h8 == myMaxDev ? GEN_2 : GEN_76;
  assign GEN_109 = 5'h9 == myMaxDev ? GEN_2 : GEN_77;
  assign GEN_110 = 5'ha == myMaxDev ? GEN_2 : GEN_78;
  assign GEN_111 = 5'hb == myMaxDev ? GEN_2 : GEN_79;
  assign GEN_112 = 5'hc == myMaxDev ? GEN_2 : GEN_80;
  assign GEN_113 = 5'hd == myMaxDev ? GEN_2 : GEN_81;
  assign GEN_114 = 5'he == myMaxDev ? GEN_2 : GEN_82;
  assign GEN_115 = 5'hf == myMaxDev ? GEN_2 : GEN_83;
  assign GEN_116 = 5'h10 == myMaxDev ? GEN_2 : GEN_84;
  assign GEN_117 = 5'h11 == myMaxDev ? GEN_2 : GEN_85;
  assign GEN_118 = 5'h12 == myMaxDev ? GEN_2 : GEN_86;
  assign GEN_119 = 5'h13 == myMaxDev ? GEN_2 : GEN_87;
  assign GEN_120 = 5'h14 == myMaxDev ? GEN_2 : GEN_88;
  assign GEN_121 = 5'h15 == myMaxDev ? GEN_2 : GEN_89;
  assign GEN_122 = 5'h16 == myMaxDev ? GEN_2 : GEN_90;
  assign GEN_123 = 5'h17 == myMaxDev ? GEN_2 : GEN_91;
  assign GEN_124 = 5'h18 == myMaxDev ? GEN_2 : GEN_92;
  assign GEN_125 = 5'h19 == myMaxDev ? GEN_2 : GEN_93;
  assign GEN_126 = 5'h1a == myMaxDev ? GEN_2 : GEN_94;
  assign GEN_127 = 5'h1b == myMaxDev ? GEN_2 : GEN_95;
  assign GEN_128 = 5'h1c == myMaxDev ? GEN_2 : GEN_96;
  assign GEN_129 = 5'h1d == myMaxDev ? GEN_2 : GEN_97;
  assign GEN_130 = 5'h1e == myMaxDev ? GEN_2 : GEN_98;
  assign GEN_131 = 5'h1f == myMaxDev ? GEN_2 : GEN_99;
  assign GEN_134 = T_1415 ? GEN_101 : GEN_69;
  assign GEN_135 = T_1415 ? GEN_102 : GEN_70;
  assign GEN_136 = T_1415 ? GEN_103 : GEN_71;
  assign GEN_137 = T_1415 ? GEN_104 : GEN_72;
  assign GEN_138 = T_1415 ? GEN_105 : GEN_73;
  assign GEN_139 = T_1415 ? GEN_106 : GEN_74;
  assign GEN_140 = T_1415 ? GEN_107 : GEN_75;
  assign GEN_141 = T_1415 ? GEN_108 : GEN_76;
  assign GEN_142 = T_1415 ? GEN_109 : GEN_77;
  assign GEN_143 = T_1415 ? GEN_110 : GEN_78;
  assign GEN_144 = T_1415 ? GEN_111 : GEN_79;
  assign GEN_145 = T_1415 ? GEN_112 : GEN_80;
  assign GEN_146 = T_1415 ? GEN_113 : GEN_81;
  assign GEN_147 = T_1415 ? GEN_114 : GEN_82;
  assign GEN_148 = T_1415 ? GEN_115 : GEN_83;
  assign GEN_149 = T_1415 ? GEN_116 : GEN_84;
  assign GEN_150 = T_1415 ? GEN_117 : GEN_85;
  assign GEN_151 = T_1415 ? GEN_118 : GEN_86;
  assign GEN_152 = T_1415 ? GEN_119 : GEN_87;
  assign GEN_153 = T_1415 ? GEN_120 : GEN_88;
  assign GEN_154 = T_1415 ? GEN_121 : GEN_89;
  assign GEN_155 = T_1415 ? GEN_122 : GEN_90;
  assign GEN_156 = T_1415 ? GEN_123 : GEN_91;
  assign GEN_157 = T_1415 ? GEN_124 : GEN_92;
  assign GEN_158 = T_1415 ? GEN_125 : GEN_93;
  assign GEN_159 = T_1415 ? GEN_126 : GEN_94;
  assign GEN_160 = T_1415 ? GEN_127 : GEN_95;
  assign GEN_161 = T_1415 ? GEN_128 : GEN_96;
  assign GEN_162 = T_1415 ? GEN_129 : GEN_97;
  assign GEN_163 = T_1415 ? GEN_130 : GEN_98;
  assign GEN_164 = T_1415 ? GEN_131 : GEN_99;
  assign T_1447 = acq_io_deq_bits_data[63:32];
  assign T_1448 = T_1447[4:0];
  assign GEN_3 = GEN_195;
  assign GEN_717 = 1'h0 == hart;
  assign GEN_718 = 5'h1 == T_1448;
  assign GEN_165 = GEN_717 & GEN_718 ? enables_0_1 : enables_0_0;
  assign GEN_720 = 5'h2 == T_1448;
  assign GEN_166 = GEN_717 & GEN_720 ? enables_0_2 : GEN_165;
  assign GEN_722 = 5'h3 == T_1448;
  assign GEN_167 = GEN_717 & GEN_722 ? enables_0_3 : GEN_166;
  assign GEN_724 = 5'h4 == T_1448;
  assign GEN_168 = GEN_717 & GEN_724 ? enables_0_4 : GEN_167;
  assign GEN_726 = 5'h5 == T_1448;
  assign GEN_169 = GEN_717 & GEN_726 ? enables_0_5 : GEN_168;
  assign GEN_728 = 5'h6 == T_1448;
  assign GEN_170 = GEN_717 & GEN_728 ? enables_0_6 : GEN_169;
  assign GEN_730 = 5'h7 == T_1448;
  assign GEN_171 = GEN_717 & GEN_730 ? enables_0_7 : GEN_170;
  assign GEN_732 = 5'h8 == T_1448;
  assign GEN_172 = GEN_717 & GEN_732 ? enables_0_8 : GEN_171;
  assign GEN_734 = 5'h9 == T_1448;
  assign GEN_173 = GEN_717 & GEN_734 ? enables_0_9 : GEN_172;
  assign GEN_736 = 5'ha == T_1448;
  assign GEN_174 = GEN_717 & GEN_736 ? enables_0_10 : GEN_173;
  assign GEN_738 = 5'hb == T_1448;
  assign GEN_175 = GEN_717 & GEN_738 ? enables_0_11 : GEN_174;
  assign GEN_740 = 5'hc == T_1448;
  assign GEN_176 = GEN_717 & GEN_740 ? enables_0_12 : GEN_175;
  assign GEN_742 = 5'hd == T_1448;
  assign GEN_177 = GEN_717 & GEN_742 ? enables_0_13 : GEN_176;
  assign GEN_744 = 5'he == T_1448;
  assign GEN_178 = GEN_717 & GEN_744 ? enables_0_14 : GEN_177;
  assign GEN_746 = 5'hf == T_1448;
  assign GEN_179 = GEN_717 & GEN_746 ? enables_0_15 : GEN_178;
  assign GEN_748 = 5'h10 == T_1448;
  assign GEN_180 = GEN_717 & GEN_748 ? enables_0_16 : GEN_179;
  assign GEN_750 = 5'h11 == T_1448;
  assign GEN_181 = GEN_717 & GEN_750 ? enables_0_17 : GEN_180;
  assign GEN_752 = 5'h12 == T_1448;
  assign GEN_182 = GEN_717 & GEN_752 ? enables_0_18 : GEN_181;
  assign GEN_754 = 5'h13 == T_1448;
  assign GEN_183 = GEN_717 & GEN_754 ? enables_0_19 : GEN_182;
  assign GEN_756 = 5'h14 == T_1448;
  assign GEN_184 = GEN_717 & GEN_756 ? enables_0_20 : GEN_183;
  assign GEN_758 = 5'h15 == T_1448;
  assign GEN_185 = GEN_717 & GEN_758 ? enables_0_21 : GEN_184;
  assign GEN_760 = 5'h16 == T_1448;
  assign GEN_186 = GEN_717 & GEN_760 ? enables_0_22 : GEN_185;
  assign GEN_762 = 5'h17 == T_1448;
  assign GEN_187 = GEN_717 & GEN_762 ? enables_0_23 : GEN_186;
  assign GEN_764 = 5'h18 == T_1448;
  assign GEN_188 = GEN_717 & GEN_764 ? enables_0_24 : GEN_187;
  assign GEN_766 = 5'h19 == T_1448;
  assign GEN_189 = GEN_717 & GEN_766 ? enables_0_25 : GEN_188;
  assign GEN_768 = 5'h1a == T_1448;
  assign GEN_190 = GEN_717 & GEN_768 ? enables_0_26 : GEN_189;
  assign GEN_770 = 5'h1b == T_1448;
  assign GEN_191 = GEN_717 & GEN_770 ? enables_0_27 : GEN_190;
  assign GEN_772 = 5'h1c == T_1448;
  assign GEN_192 = GEN_717 & GEN_772 ? enables_0_28 : GEN_191;
  assign GEN_774 = 5'h1d == T_1448;
  assign GEN_193 = GEN_717 & GEN_774 ? enables_0_29 : GEN_192;
  assign GEN_776 = 5'h1e == T_1448;
  assign GEN_194 = GEN_717 & GEN_776 ? enables_0_30 : GEN_193;
  assign GEN_778 = 5'h1f == T_1448;
  assign GEN_195 = GEN_717 & GEN_778 ? enables_0_31 : GEN_194;
  assign T_1450 = T_1448 - 5'h1;
  assign T_1451 = T_1450[4:0];
  assign GEN_4 = 1'h1;
  assign GEN_196 = 5'h0 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_197 = 5'h1 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_198 = 5'h2 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_199 = 5'h3 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_200 = 5'h4 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_201 = 5'h5 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_202 = 5'h6 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_203 = 5'h7 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_204 = 5'h8 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_205 = 5'h9 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_206 = 5'ha == T_1451 ? GEN_4 : 1'h0;
  assign GEN_207 = 5'hb == T_1451 ? GEN_4 : 1'h0;
  assign GEN_208 = 5'hc == T_1451 ? GEN_4 : 1'h0;
  assign GEN_209 = 5'hd == T_1451 ? GEN_4 : 1'h0;
  assign GEN_210 = 5'he == T_1451 ? GEN_4 : 1'h0;
  assign GEN_211 = 5'hf == T_1451 ? GEN_4 : 1'h0;
  assign GEN_212 = 5'h10 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_213 = 5'h11 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_214 = 5'h12 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_215 = 5'h13 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_216 = 5'h14 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_217 = 5'h15 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_218 = 5'h16 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_219 = 5'h17 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_220 = 5'h18 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_221 = 5'h19 == T_1451 ? GEN_4 : 1'h0;
  assign GEN_222 = 5'h1a == T_1451 ? GEN_4 : 1'h0;
  assign GEN_223 = 5'h1b == T_1451 ? GEN_4 : 1'h0;
  assign GEN_224 = 5'h1c == T_1451 ? GEN_4 : 1'h0;
  assign GEN_225 = 5'h1d == T_1451 ? GEN_4 : 1'h0;
  assign GEN_226 = 5'h1e == T_1451 ? GEN_4 : 1'h0;
  assign GEN_228 = GEN_3 ? GEN_196 : 1'h0;
  assign GEN_229 = GEN_3 ? GEN_197 : 1'h0;
  assign GEN_230 = GEN_3 ? GEN_198 : 1'h0;
  assign GEN_231 = GEN_3 ? GEN_199 : 1'h0;
  assign GEN_232 = GEN_3 ? GEN_200 : 1'h0;
  assign GEN_233 = GEN_3 ? GEN_201 : 1'h0;
  assign GEN_234 = GEN_3 ? GEN_202 : 1'h0;
  assign GEN_235 = GEN_3 ? GEN_203 : 1'h0;
  assign GEN_236 = GEN_3 ? GEN_204 : 1'h0;
  assign GEN_237 = GEN_3 ? GEN_205 : 1'h0;
  assign GEN_238 = GEN_3 ? GEN_206 : 1'h0;
  assign GEN_239 = GEN_3 ? GEN_207 : 1'h0;
  assign GEN_240 = GEN_3 ? GEN_208 : 1'h0;
  assign GEN_241 = GEN_3 ? GEN_209 : 1'h0;
  assign GEN_242 = GEN_3 ? GEN_210 : 1'h0;
  assign GEN_243 = GEN_3 ? GEN_211 : 1'h0;
  assign GEN_244 = GEN_3 ? GEN_212 : 1'h0;
  assign GEN_245 = GEN_3 ? GEN_213 : 1'h0;
  assign GEN_246 = GEN_3 ? GEN_214 : 1'h0;
  assign GEN_247 = GEN_3 ? GEN_215 : 1'h0;
  assign GEN_248 = GEN_3 ? GEN_216 : 1'h0;
  assign GEN_249 = GEN_3 ? GEN_217 : 1'h0;
  assign GEN_250 = GEN_3 ? GEN_218 : 1'h0;
  assign GEN_251 = GEN_3 ? GEN_219 : 1'h0;
  assign GEN_252 = GEN_3 ? GEN_220 : 1'h0;
  assign GEN_253 = GEN_3 ? GEN_221 : 1'h0;
  assign GEN_254 = GEN_3 ? GEN_222 : 1'h0;
  assign GEN_255 = GEN_3 ? GEN_223 : 1'h0;
  assign GEN_256 = GEN_3 ? GEN_224 : 1'h0;
  assign GEN_257 = GEN_3 ? GEN_225 : 1'h0;
  assign GEN_258 = GEN_3 ? GEN_226 : 1'h0;
  assign GEN_261 = T_1283 ? GEN_228 : 1'h0;
  assign GEN_262 = T_1283 ? GEN_229 : 1'h0;
  assign GEN_263 = T_1283 ? GEN_230 : 1'h0;
  assign GEN_264 = T_1283 ? GEN_231 : 1'h0;
  assign GEN_265 = T_1283 ? GEN_232 : 1'h0;
  assign GEN_266 = T_1283 ? GEN_233 : 1'h0;
  assign GEN_267 = T_1283 ? GEN_234 : 1'h0;
  assign GEN_268 = T_1283 ? GEN_235 : 1'h0;
  assign GEN_269 = T_1283 ? GEN_236 : 1'h0;
  assign GEN_270 = T_1283 ? GEN_237 : 1'h0;
  assign GEN_271 = T_1283 ? GEN_238 : 1'h0;
  assign GEN_272 = T_1283 ? GEN_239 : 1'h0;
  assign GEN_273 = T_1283 ? GEN_240 : 1'h0;
  assign GEN_274 = T_1283 ? GEN_241 : 1'h0;
  assign GEN_275 = T_1283 ? GEN_242 : 1'h0;
  assign GEN_276 = T_1283 ? GEN_243 : 1'h0;
  assign GEN_277 = T_1283 ? GEN_244 : 1'h0;
  assign GEN_278 = T_1283 ? GEN_245 : 1'h0;
  assign GEN_279 = T_1283 ? GEN_246 : 1'h0;
  assign GEN_280 = T_1283 ? GEN_247 : 1'h0;
  assign GEN_281 = T_1283 ? GEN_248 : 1'h0;
  assign GEN_282 = T_1283 ? GEN_249 : 1'h0;
  assign GEN_283 = T_1283 ? GEN_250 : 1'h0;
  assign GEN_284 = T_1283 ? GEN_251 : 1'h0;
  assign GEN_285 = T_1283 ? GEN_252 : 1'h0;
  assign GEN_286 = T_1283 ? GEN_253 : 1'h0;
  assign GEN_287 = T_1283 ? GEN_254 : 1'h0;
  assign GEN_288 = T_1283 ? GEN_255 : 1'h0;
  assign GEN_289 = T_1283 ? GEN_256 : 1'h0;
  assign GEN_290 = T_1283 ? GEN_257 : 1'h0;
  assign GEN_291 = T_1283 ? GEN_258 : 1'h0;
  assign GEN_294 = write ? GEN_261 : 1'h0;
  assign GEN_295 = write ? GEN_262 : 1'h0;
  assign GEN_296 = write ? GEN_263 : 1'h0;
  assign GEN_297 = write ? GEN_264 : 1'h0;
  assign GEN_298 = write ? GEN_265 : 1'h0;
  assign GEN_299 = write ? GEN_266 : 1'h0;
  assign GEN_300 = write ? GEN_267 : 1'h0;
  assign GEN_301 = write ? GEN_268 : 1'h0;
  assign GEN_302 = write ? GEN_269 : 1'h0;
  assign GEN_303 = write ? GEN_270 : 1'h0;
  assign GEN_304 = write ? GEN_271 : 1'h0;
  assign GEN_305 = write ? GEN_272 : 1'h0;
  assign GEN_306 = write ? GEN_273 : 1'h0;
  assign GEN_307 = write ? GEN_274 : 1'h0;
  assign GEN_308 = write ? GEN_275 : 1'h0;
  assign GEN_309 = write ? GEN_276 : 1'h0;
  assign GEN_310 = write ? GEN_277 : 1'h0;
  assign GEN_311 = write ? GEN_278 : 1'h0;
  assign GEN_312 = write ? GEN_279 : 1'h0;
  assign GEN_313 = write ? GEN_280 : 1'h0;
  assign GEN_314 = write ? GEN_281 : 1'h0;
  assign GEN_315 = write ? GEN_282 : 1'h0;
  assign GEN_316 = write ? GEN_283 : 1'h0;
  assign GEN_317 = write ? GEN_284 : 1'h0;
  assign GEN_318 = write ? GEN_285 : 1'h0;
  assign GEN_319 = write ? GEN_286 : 1'h0;
  assign GEN_320 = write ? GEN_287 : 1'h0;
  assign GEN_321 = write ? GEN_288 : 1'h0;
  assign GEN_322 = write ? GEN_289 : 1'h0;
  assign GEN_323 = write ? GEN_290 : 1'h0;
  assign GEN_324 = write ? GEN_291 : 1'h0;
  assign GEN_326 = T_1406 ? {{27'd0}, T_1413} : 64'h0;
  assign GEN_329 = T_1406 ? GEN_134 : GEN_69;
  assign GEN_330 = T_1406 ? GEN_135 : GEN_70;
  assign GEN_331 = T_1406 ? GEN_136 : GEN_71;
  assign GEN_332 = T_1406 ? GEN_137 : GEN_72;
  assign GEN_333 = T_1406 ? GEN_138 : GEN_73;
  assign GEN_334 = T_1406 ? GEN_139 : GEN_74;
  assign GEN_335 = T_1406 ? GEN_140 : GEN_75;
  assign GEN_336 = T_1406 ? GEN_141 : GEN_76;
  assign GEN_337 = T_1406 ? GEN_142 : GEN_77;
  assign GEN_338 = T_1406 ? GEN_143 : GEN_78;
  assign GEN_339 = T_1406 ? GEN_144 : GEN_79;
  assign GEN_340 = T_1406 ? GEN_145 : GEN_80;
  assign GEN_341 = T_1406 ? GEN_146 : GEN_81;
  assign GEN_342 = T_1406 ? GEN_147 : GEN_82;
  assign GEN_343 = T_1406 ? GEN_148 : GEN_83;
  assign GEN_344 = T_1406 ? GEN_149 : GEN_84;
  assign GEN_345 = T_1406 ? GEN_150 : GEN_85;
  assign GEN_346 = T_1406 ? GEN_151 : GEN_86;
  assign GEN_347 = T_1406 ? GEN_152 : GEN_87;
  assign GEN_348 = T_1406 ? GEN_153 : GEN_88;
  assign GEN_349 = T_1406 ? GEN_154 : GEN_89;
  assign GEN_350 = T_1406 ? GEN_155 : GEN_90;
  assign GEN_351 = T_1406 ? GEN_156 : GEN_91;
  assign GEN_352 = T_1406 ? GEN_157 : GEN_92;
  assign GEN_353 = T_1406 ? GEN_158 : GEN_93;
  assign GEN_354 = T_1406 ? GEN_159 : GEN_94;
  assign GEN_355 = T_1406 ? GEN_160 : GEN_95;
  assign GEN_356 = T_1406 ? GEN_161 : GEN_96;
  assign GEN_357 = T_1406 ? GEN_162 : GEN_97;
  assign GEN_358 = T_1406 ? GEN_163 : GEN_98;
  assign GEN_359 = T_1406 ? GEN_164 : GEN_99;
  assign GEN_362 = T_1406 ? GEN_294 : 1'h0;
  assign GEN_363 = T_1406 ? GEN_295 : 1'h0;
  assign GEN_364 = T_1406 ? GEN_296 : 1'h0;
  assign GEN_365 = T_1406 ? GEN_297 : 1'h0;
  assign GEN_366 = T_1406 ? GEN_298 : 1'h0;
  assign GEN_367 = T_1406 ? GEN_299 : 1'h0;
  assign GEN_368 = T_1406 ? GEN_300 : 1'h0;
  assign GEN_369 = T_1406 ? GEN_301 : 1'h0;
  assign GEN_370 = T_1406 ? GEN_302 : 1'h0;
  assign GEN_371 = T_1406 ? GEN_303 : 1'h0;
  assign GEN_372 = T_1406 ? GEN_304 : 1'h0;
  assign GEN_373 = T_1406 ? GEN_305 : 1'h0;
  assign GEN_374 = T_1406 ? GEN_306 : 1'h0;
  assign GEN_375 = T_1406 ? GEN_307 : 1'h0;
  assign GEN_376 = T_1406 ? GEN_308 : 1'h0;
  assign GEN_377 = T_1406 ? GEN_309 : 1'h0;
  assign GEN_378 = T_1406 ? GEN_310 : 1'h0;
  assign GEN_379 = T_1406 ? GEN_311 : 1'h0;
  assign GEN_380 = T_1406 ? GEN_312 : 1'h0;
  assign GEN_381 = T_1406 ? GEN_313 : 1'h0;
  assign GEN_382 = T_1406 ? GEN_314 : 1'h0;
  assign GEN_383 = T_1406 ? GEN_315 : 1'h0;
  assign GEN_384 = T_1406 ? GEN_316 : 1'h0;
  assign GEN_385 = T_1406 ? GEN_317 : 1'h0;
  assign GEN_386 = T_1406 ? GEN_318 : 1'h0;
  assign GEN_387 = T_1406 ? GEN_319 : 1'h0;
  assign GEN_388 = T_1406 ? GEN_320 : 1'h0;
  assign GEN_389 = T_1406 ? GEN_321 : 1'h0;
  assign GEN_390 = T_1406 ? GEN_322 : 1'h0;
  assign GEN_391 = T_1406 ? GEN_323 : 1'h0;
  assign GEN_392 = T_1406 ? GEN_324 : 1'h0;
  assign T_1459 = addr >= 26'h2000;
  assign T_1461 = T_1406 == 1'h0;
  assign T_1462 = T_1461 & T_1459;
  assign GEN_5 = enables_0_1;
  assign GEN_6 = enables_0_0;
  assign T_1467 = {GEN_5,GEN_6};
  assign GEN_7 = enables_0_3;
  assign GEN_8 = enables_0_2;
  assign T_1468 = {GEN_7,GEN_8};
  assign T_1469 = {T_1468,T_1467};
  assign GEN_9 = enables_0_5;
  assign GEN_10 = enables_0_4;
  assign T_1470 = {GEN_9,GEN_10};
  assign GEN_11 = enables_0_7;
  assign GEN_12 = enables_0_6;
  assign T_1471 = {GEN_11,GEN_12};
  assign T_1472 = {T_1471,T_1470};
  assign T_1473 = {T_1472,T_1469};
  assign GEN_13 = enables_0_9;
  assign GEN_14 = enables_0_8;
  assign T_1474 = {GEN_13,GEN_14};
  assign GEN_15 = enables_0_11;
  assign GEN_16 = enables_0_10;
  assign T_1475 = {GEN_15,GEN_16};
  assign T_1476 = {T_1475,T_1474};
  assign GEN_17 = enables_0_13;
  assign GEN_18 = enables_0_12;
  assign T_1477 = {GEN_17,GEN_18};
  assign GEN_19 = enables_0_15;
  assign GEN_20 = enables_0_14;
  assign T_1478 = {GEN_19,GEN_20};
  assign T_1479 = {T_1478,T_1477};
  assign T_1480 = {T_1479,T_1476};
  assign T_1481 = {T_1480,T_1473};
  assign GEN_21 = enables_0_17;
  assign GEN_22 = enables_0_16;
  assign T_1482 = {GEN_21,GEN_22};
  assign GEN_23 = enables_0_19;
  assign GEN_24 = enables_0_18;
  assign T_1483 = {GEN_23,GEN_24};
  assign T_1484 = {T_1483,T_1482};
  assign GEN_25 = enables_0_21;
  assign GEN_26 = enables_0_20;
  assign T_1485 = {GEN_25,GEN_26};
  assign GEN_27 = enables_0_23;
  assign GEN_28 = enables_0_22;
  assign T_1486 = {GEN_27,GEN_28};
  assign T_1487 = {T_1486,T_1485};
  assign T_1488 = {T_1487,T_1484};
  assign GEN_29 = enables_0_25;
  assign GEN_30 = enables_0_24;
  assign T_1489 = {GEN_29,GEN_30};
  assign GEN_31 = enables_0_27;
  assign GEN_32 = enables_0_26;
  assign T_1490 = {GEN_31,GEN_32};
  assign T_1491 = {T_1490,T_1489};
  assign GEN_33 = enables_0_29;
  assign GEN_34 = enables_0_28;
  assign T_1492 = {GEN_33,GEN_34};
  assign GEN_35 = enables_0_31;
  assign GEN_36 = enables_0_30;
  assign T_1493 = {GEN_35,GEN_36};
  assign T_1494 = {T_1493,T_1492};
  assign T_1495 = {T_1494,T_1491};
  assign T_1496 = {T_1495,T_1488};
  assign T_1497 = {T_1496,T_1481};
  assign T_1501 = masked_wdata[0];
  assign GEN_37 = T_1501;
  assign T_1505 = masked_wdata[1];
  assign GEN_38 = T_1505;
  assign GEN_398 = write ? GEN_38 : enables_0_1;
  assign T_1509 = masked_wdata[2];
  assign GEN_39 = T_1509;
  assign GEN_401 = write ? GEN_39 : enables_0_2;
  assign T_1513 = masked_wdata[3];
  assign GEN_40 = T_1513;
  assign GEN_404 = write ? GEN_40 : enables_0_3;
  assign T_1517 = masked_wdata[4];
  assign GEN_41 = T_1517;
  assign GEN_407 = write ? GEN_41 : enables_0_4;
  assign T_1521 = masked_wdata[5];
  assign GEN_42 = T_1521;
  assign GEN_410 = write ? GEN_42 : enables_0_5;
  assign T_1525 = masked_wdata[6];
  assign GEN_43 = T_1525;
  assign GEN_413 = write ? GEN_43 : enables_0_6;
  assign T_1529 = masked_wdata[7];
  assign GEN_44 = T_1529;
  assign GEN_416 = write ? GEN_44 : enables_0_7;
  assign T_1533 = masked_wdata[8];
  assign GEN_45 = T_1533;
  assign GEN_419 = write ? GEN_45 : enables_0_8;
  assign T_1537 = masked_wdata[9];
  assign GEN_46 = T_1537;
  assign GEN_422 = write ? GEN_46 : enables_0_9;
  assign T_1541 = masked_wdata[10];
  assign GEN_47 = T_1541;
  assign GEN_425 = write ? GEN_47 : enables_0_10;
  assign T_1545 = masked_wdata[11];
  assign GEN_48 = T_1545;
  assign GEN_428 = write ? GEN_48 : enables_0_11;
  assign T_1549 = masked_wdata[12];
  assign GEN_49 = T_1549;
  assign GEN_431 = write ? GEN_49 : enables_0_12;
  assign T_1553 = masked_wdata[13];
  assign GEN_50 = T_1553;
  assign GEN_434 = write ? GEN_50 : enables_0_13;
  assign T_1557 = masked_wdata[14];
  assign GEN_51 = T_1557;
  assign GEN_437 = write ? GEN_51 : enables_0_14;
  assign T_1561 = masked_wdata[15];
  assign GEN_52 = T_1561;
  assign GEN_440 = write ? GEN_52 : enables_0_15;
  assign T_1565 = masked_wdata[16];
  assign GEN_53 = T_1565;
  assign GEN_443 = write ? GEN_53 : enables_0_16;
  assign T_1569 = masked_wdata[17];
  assign GEN_54 = T_1569;
  assign GEN_446 = write ? GEN_54 : enables_0_17;
  assign T_1573 = masked_wdata[18];
  assign GEN_55 = T_1573;
  assign GEN_449 = write ? GEN_55 : enables_0_18;
  assign T_1577 = masked_wdata[19];
  assign GEN_56 = T_1577;
  assign GEN_452 = write ? GEN_56 : enables_0_19;
  assign T_1581 = masked_wdata[20];
  assign GEN_57 = T_1581;
  assign GEN_455 = write ? GEN_57 : enables_0_20;
  assign T_1585 = masked_wdata[21];
  assign GEN_58 = T_1585;
  assign GEN_458 = write ? GEN_58 : enables_0_21;
  assign T_1589 = masked_wdata[22];
  assign GEN_59 = T_1589;
  assign GEN_461 = write ? GEN_59 : enables_0_22;
  assign T_1593 = masked_wdata[23];
  assign GEN_60 = T_1593;
  assign GEN_464 = write ? GEN_60 : enables_0_23;
  assign T_1597 = masked_wdata[24];
  assign GEN_61 = T_1597;
  assign GEN_467 = write ? GEN_61 : enables_0_24;
  assign T_1601 = masked_wdata[25];
  assign GEN_62 = T_1601;
  assign GEN_470 = write ? GEN_62 : enables_0_25;
  assign T_1605 = masked_wdata[26];
  assign GEN_63 = T_1605;
  assign GEN_473 = write ? GEN_63 : enables_0_26;
  assign T_1609 = masked_wdata[27];
  assign GEN_64 = T_1609;
  assign GEN_476 = write ? GEN_64 : enables_0_27;
  assign T_1613 = masked_wdata[28];
  assign GEN_65 = T_1613;
  assign GEN_479 = write ? GEN_65 : enables_0_28;
  assign T_1617 = masked_wdata[29];
  assign GEN_66 = T_1617;
  assign GEN_482 = write ? GEN_66 : enables_0_29;
  assign T_1621 = masked_wdata[30];
  assign GEN_67 = T_1621;
  assign GEN_485 = write ? GEN_67 : enables_0_30;
  assign T_1625 = masked_wdata[31];
  assign GEN_68 = T_1625;
  assign GEN_488 = write ? GEN_68 : enables_0_31;
  assign GEN_521 = {{32'd0}, T_1497};
  assign GEN_619 = T_1462 ? GEN_521 : GEN_326;
  assign GEN_623 = T_1462 ? GEN_398 : enables_0_1;
  assign GEN_625 = T_1462 ? GEN_401 : enables_0_2;
  assign GEN_627 = T_1462 ? GEN_404 : enables_0_3;
  assign GEN_629 = T_1462 ? GEN_407 : enables_0_4;
  assign GEN_631 = T_1462 ? GEN_410 : enables_0_5;
  assign GEN_633 = T_1462 ? GEN_413 : enables_0_6;
  assign GEN_635 = T_1462 ? GEN_416 : enables_0_7;
  assign GEN_637 = T_1462 ? GEN_419 : enables_0_8;
  assign GEN_639 = T_1462 ? GEN_422 : enables_0_9;
  assign GEN_641 = T_1462 ? GEN_425 : enables_0_10;
  assign GEN_643 = T_1462 ? GEN_428 : enables_0_11;
  assign GEN_645 = T_1462 ? GEN_431 : enables_0_12;
  assign GEN_647 = T_1462 ? GEN_434 : enables_0_13;
  assign GEN_649 = T_1462 ? GEN_437 : enables_0_14;
  assign GEN_651 = T_1462 ? GEN_440 : enables_0_15;
  assign GEN_653 = T_1462 ? GEN_443 : enables_0_16;
  assign GEN_655 = T_1462 ? GEN_446 : enables_0_17;
  assign GEN_657 = T_1462 ? GEN_449 : enables_0_18;
  assign GEN_659 = T_1462 ? GEN_452 : enables_0_19;
  assign GEN_661 = T_1462 ? GEN_455 : enables_0_20;
  assign GEN_663 = T_1462 ? GEN_458 : enables_0_21;
  assign GEN_665 = T_1462 ? GEN_461 : enables_0_22;
  assign GEN_667 = T_1462 ? GEN_464 : enables_0_23;
  assign GEN_669 = T_1462 ? GEN_467 : enables_0_24;
  assign GEN_671 = T_1462 ? GEN_470 : enables_0_25;
  assign GEN_673 = T_1462 ? GEN_473 : enables_0_26;
  assign GEN_675 = T_1462 ? GEN_476 : enables_0_27;
  assign GEN_677 = T_1462 ? GEN_479 : enables_0_28;
  assign GEN_679 = T_1462 ? GEN_482 : enables_0_29;
  assign GEN_681 = T_1462 ? GEN_485 : enables_0_30;
  assign GEN_683 = T_1462 ? GEN_488 : enables_0_31;
  assign T_1627 = addr >= 26'h1000;
  assign T_1631 = T_1459 == 1'h0;
  assign T_1632 = T_1461 & T_1631;
  assign T_1633 = T_1632 & T_1627;
  assign T_1634 = addr[4:3];
  assign T_1635 = {pending_1,pending_0};
  assign T_1636 = {pending_3,pending_2};
  assign T_1637 = {T_1636,T_1635};
  assign T_1638 = {pending_5,pending_4};
  assign T_1639 = {pending_7,pending_6};
  assign T_1640 = {T_1639,T_1638};
  assign T_1641 = {T_1640,T_1637};
  assign T_1642 = {pending_9,pending_8};
  assign T_1643 = {pending_11,pending_10};
  assign T_1644 = {T_1643,T_1642};
  assign T_1645 = {pending_13,pending_12};
  assign T_1646 = {pending_15,pending_14};
  assign T_1647 = {T_1646,T_1645};
  assign T_1648 = {T_1647,T_1644};
  assign T_1649 = {T_1648,T_1641};
  assign T_1650 = {pending_17,pending_16};
  assign T_1651 = {pending_19,pending_18};
  assign T_1652 = {T_1651,T_1650};
  assign T_1653 = {pending_21,pending_20};
  assign T_1654 = {pending_23,pending_22};
  assign T_1655 = {T_1654,T_1653};
  assign T_1656 = {T_1655,T_1652};
  assign T_1657 = {pending_25,pending_24};
  assign T_1658 = {pending_27,pending_26};
  assign T_1659 = {T_1658,T_1657};
  assign T_1660 = {pending_29,pending_28};
  assign T_1661 = {pending_31,pending_30};
  assign T_1662 = {T_1661,T_1660};
  assign T_1663 = {T_1662,T_1659};
  assign T_1664 = {T_1663,T_1656};
  assign T_1665 = {T_1664,T_1649};
  assign GEN_779 = {{5'd0}, T_1634};
  assign T_1667 = GEN_779 * 7'h40;
  assign T_1668 = T_1665 >> T_1667;
  assign GEN_684 = T_1633 ? {{32'd0}, T_1668} : GEN_619;
  assign T_1675 = T_1627 == 1'h0;
  assign T_1676 = T_1632 & T_1675;
  assign T_1677 = addr[6:3];
  assign T_1679 = T_1677 == 4'h0;
  assign T_1681 = {31'h0,priority_0};
  assign T_1683 = {31'h0,priority_1};
  assign T_1684 = {T_1683,T_1681};
  assign GEN_685 = T_1679 ? T_1684 : GEN_684;
  assign T_1686 = T_1677 == 4'h1;
  assign T_1688 = {31'h0,priority_2};
  assign T_1690 = {31'h0,priority_3};
  assign T_1691 = {T_1690,T_1688};
  assign GEN_686 = T_1686 ? T_1691 : GEN_685;
  assign T_1693 = T_1677 == 4'h2;
  assign T_1695 = {31'h0,priority_4};
  assign T_1697 = {31'h0,priority_5};
  assign T_1698 = {T_1697,T_1695};
  assign GEN_687 = T_1693 ? T_1698 : GEN_686;
  assign T_1700 = T_1677 == 4'h3;
  assign T_1702 = {31'h0,priority_6};
  assign T_1704 = {31'h0,priority_7};
  assign T_1705 = {T_1704,T_1702};
  assign GEN_688 = T_1700 ? T_1705 : GEN_687;
  assign T_1707 = T_1677 == 4'h4;
  assign T_1709 = {31'h0,priority_8};
  assign T_1711 = {31'h0,priority_9};
  assign T_1712 = {T_1711,T_1709};
  assign GEN_689 = T_1707 ? T_1712 : GEN_688;
  assign T_1714 = T_1677 == 4'h5;
  assign T_1716 = {31'h0,priority_10};
  assign T_1718 = {31'h0,priority_11};
  assign T_1719 = {T_1718,T_1716};
  assign GEN_690 = T_1714 ? T_1719 : GEN_689;
  assign T_1721 = T_1677 == 4'h6;
  assign T_1723 = {31'h0,priority_12};
  assign T_1725 = {31'h0,priority_13};
  assign T_1726 = {T_1725,T_1723};
  assign GEN_691 = T_1721 ? T_1726 : GEN_690;
  assign T_1728 = T_1677 == 4'h7;
  assign T_1730 = {31'h0,priority_14};
  assign T_1732 = {31'h0,priority_15};
  assign T_1733 = {T_1732,T_1730};
  assign GEN_692 = T_1728 ? T_1733 : GEN_691;
  assign T_1735 = T_1677 == 4'h8;
  assign T_1737 = {31'h0,priority_16};
  assign T_1739 = {31'h0,priority_17};
  assign T_1740 = {T_1739,T_1737};
  assign GEN_693 = T_1735 ? T_1740 : GEN_692;
  assign T_1742 = T_1677 == 4'h9;
  assign T_1744 = {31'h0,priority_18};
  assign T_1746 = {31'h0,priority_19};
  assign T_1747 = {T_1746,T_1744};
  assign GEN_694 = T_1742 ? T_1747 : GEN_693;
  assign T_1749 = T_1677 == 4'ha;
  assign T_1751 = {31'h0,priority_20};
  assign T_1753 = {31'h0,priority_21};
  assign T_1754 = {T_1753,T_1751};
  assign GEN_695 = T_1749 ? T_1754 : GEN_694;
  assign T_1756 = T_1677 == 4'hb;
  assign T_1758 = {31'h0,priority_22};
  assign T_1760 = {31'h0,priority_23};
  assign T_1761 = {T_1760,T_1758};
  assign GEN_696 = T_1756 ? T_1761 : GEN_695;
  assign T_1763 = T_1677 == 4'hc;
  assign T_1765 = {31'h0,priority_24};
  assign T_1767 = {31'h0,priority_25};
  assign T_1768 = {T_1767,T_1765};
  assign GEN_697 = T_1763 ? T_1768 : GEN_696;
  assign T_1770 = T_1677 == 4'hd;
  assign T_1772 = {31'h0,priority_26};
  assign T_1774 = {31'h0,priority_27};
  assign T_1775 = {T_1774,T_1772};
  assign GEN_698 = T_1770 ? T_1775 : GEN_697;
  assign T_1777 = T_1677 == 4'he;
  assign T_1779 = {31'h0,priority_28};
  assign T_1781 = {31'h0,priority_29};
  assign T_1782 = {T_1781,T_1779};
  assign GEN_699 = T_1777 ? T_1782 : GEN_698;
  assign T_1784 = T_1677 == 4'hf;
  assign T_1786 = {31'h0,priority_30};
  assign T_1788 = {31'h0,priority_31};
  assign T_1789 = {T_1788,T_1786};
  assign GEN_700 = T_1784 ? T_1789 : GEN_699;
  assign GEN_701 = T_1676 ? GEN_700 : GEN_684;
  assign T_1809 = 3'h6 == acq_io_deq_bits_a_type;
  assign T_1810 = T_1809 ? 3'h1 : 3'h3;
  assign T_1811 = 3'h5 == acq_io_deq_bits_a_type;
  assign T_1812 = T_1811 ? 3'h1 : T_1810;
  assign T_1813 = 3'h4 == acq_io_deq_bits_a_type;
  assign T_1814 = T_1813 ? 3'h4 : T_1812;
  assign T_1815 = 3'h3 == acq_io_deq_bits_a_type;
  assign T_1816 = T_1815 ? 3'h3 : T_1814;
  assign T_1817 = 3'h2 == acq_io_deq_bits_a_type;
  assign T_1818 = T_1817 ? 3'h3 : T_1816;
  assign T_1819 = 3'h1 == acq_io_deq_bits_a_type;
  assign T_1820 = T_1819 ? 3'h5 : T_1818;
  assign T_1821 = 3'h0 == acq_io_deq_bits_a_type;
  assign T_1822 = T_1821 ? 3'h4 : T_1820;
  assign T_1847_addr_beat = 3'h0;
  assign T_1847_client_xact_id = acq_io_deq_bits_client_xact_id;
  assign T_1847_manager_xact_id = 1'h0;
  assign T_1847_is_builtin_type = 1'h1;
  assign T_1847_g_type = {{1'd0}, T_1822};
  assign T_1847_data = rdata;
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002;
    `endif
  `ifdef RANDOMIZE
  GEN_100 = {1{$random}};
  pending_0 = GEN_100[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_132 = {1{$random}};
  pending_1 = GEN_132[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_133 = {1{$random}};
  pending_2 = GEN_133[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_227 = {1{$random}};
  pending_3 = GEN_227[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_259 = {1{$random}};
  pending_4 = GEN_259[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_260 = {1{$random}};
  pending_5 = GEN_260[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_292 = {1{$random}};
  pending_6 = GEN_292[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_293 = {1{$random}};
  pending_7 = GEN_293[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_325 = {1{$random}};
  pending_8 = GEN_325[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_327 = {1{$random}};
  pending_9 = GEN_327[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_328 = {1{$random}};
  pending_10 = GEN_328[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_360 = {1{$random}};
  pending_11 = GEN_360[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_361 = {1{$random}};
  pending_12 = GEN_361[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_393 = {1{$random}};
  pending_13 = GEN_393[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_394 = {1{$random}};
  pending_14 = GEN_394[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_395 = {1{$random}};
  pending_15 = GEN_395[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_396 = {1{$random}};
  pending_16 = GEN_396[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_397 = {1{$random}};
  pending_17 = GEN_397[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_399 = {1{$random}};
  pending_18 = GEN_399[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_400 = {1{$random}};
  pending_19 = GEN_400[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_402 = {1{$random}};
  pending_20 = GEN_402[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_403 = {1{$random}};
  pending_21 = GEN_403[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_405 = {1{$random}};
  pending_22 = GEN_405[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_406 = {1{$random}};
  pending_23 = GEN_406[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_408 = {1{$random}};
  pending_24 = GEN_408[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_409 = {1{$random}};
  pending_25 = GEN_409[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_411 = {1{$random}};
  pending_26 = GEN_411[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_412 = {1{$random}};
  pending_27 = GEN_412[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_414 = {1{$random}};
  pending_28 = GEN_414[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_415 = {1{$random}};
  pending_29 = GEN_415[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_417 = {1{$random}};
  pending_30 = GEN_417[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_418 = {1{$random}};
  pending_31 = GEN_418[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_420 = {1{$random}};
  enables_0_0 = GEN_420[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_421 = {1{$random}};
  enables_0_1 = GEN_421[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_423 = {1{$random}};
  enables_0_2 = GEN_423[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_424 = {1{$random}};
  enables_0_3 = GEN_424[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_426 = {1{$random}};
  enables_0_4 = GEN_426[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_427 = {1{$random}};
  enables_0_5 = GEN_427[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_429 = {1{$random}};
  enables_0_6 = GEN_429[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_430 = {1{$random}};
  enables_0_7 = GEN_430[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_432 = {1{$random}};
  enables_0_8 = GEN_432[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_433 = {1{$random}};
  enables_0_9 = GEN_433[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_435 = {1{$random}};
  enables_0_10 = GEN_435[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_436 = {1{$random}};
  enables_0_11 = GEN_436[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_438 = {1{$random}};
  enables_0_12 = GEN_438[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_439 = {1{$random}};
  enables_0_13 = GEN_439[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_441 = {1{$random}};
  enables_0_14 = GEN_441[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_442 = {1{$random}};
  enables_0_15 = GEN_442[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_444 = {1{$random}};
  enables_0_16 = GEN_444[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_445 = {1{$random}};
  enables_0_17 = GEN_445[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_447 = {1{$random}};
  enables_0_18 = GEN_447[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_448 = {1{$random}};
  enables_0_19 = GEN_448[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_450 = {1{$random}};
  enables_0_20 = GEN_450[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_451 = {1{$random}};
  enables_0_21 = GEN_451[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_453 = {1{$random}};
  enables_0_22 = GEN_453[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_454 = {1{$random}};
  enables_0_23 = GEN_454[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_456 = {1{$random}};
  enables_0_24 = GEN_456[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_457 = {1{$random}};
  enables_0_25 = GEN_457[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_459 = {1{$random}};
  enables_0_26 = GEN_459[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_460 = {1{$random}};
  enables_0_27 = GEN_460[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_462 = {1{$random}};
  enables_0_28 = GEN_462[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_463 = {1{$random}};
  enables_0_29 = GEN_463[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_465 = {1{$random}};
  enables_0_30 = GEN_465[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_466 = {1{$random}};
  enables_0_31 = GEN_466[0:0];
  `endif
  `ifdef RANDOMIZE
  GEN_468 = {1{$random}};
  T_1182 = GEN_468[4:0];
  `endif
  `ifdef RANDOMIZE
  GEN_469 = {1{$random}};
  T_1183 = GEN_469[1:0];
  `endif
  end
`endif
  always @(posedge clk) begin
    if(reset) begin
      pending_0 <= T_733_0;
    end else begin
      pending_0 <= 1'h0;
    end
    if(reset) begin
      pending_1 <= T_733_1;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h1 == myMaxDev) begin
            pending_1 <= GEN_2;
          end else begin
            if(io_devices_0_valid) begin
              pending_1 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_0_valid) begin
            pending_1 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_0_valid) begin
          pending_1 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_2 <= T_733_2;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h2 == myMaxDev) begin
            pending_2 <= GEN_2;
          end else begin
            if(io_devices_1_valid) begin
              pending_2 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_1_valid) begin
            pending_2 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_1_valid) begin
          pending_2 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_3 <= T_733_3;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h3 == myMaxDev) begin
            pending_3 <= GEN_2;
          end else begin
            if(io_devices_2_valid) begin
              pending_3 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_2_valid) begin
            pending_3 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_2_valid) begin
          pending_3 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_4 <= T_733_4;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h4 == myMaxDev) begin
            pending_4 <= GEN_2;
          end else begin
            if(io_devices_3_valid) begin
              pending_4 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_3_valid) begin
            pending_4 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_3_valid) begin
          pending_4 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_5 <= T_733_5;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h5 == myMaxDev) begin
            pending_5 <= GEN_2;
          end else begin
            if(io_devices_4_valid) begin
              pending_5 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_4_valid) begin
            pending_5 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_4_valid) begin
          pending_5 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_6 <= T_733_6;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h6 == myMaxDev) begin
            pending_6 <= GEN_2;
          end else begin
            if(io_devices_5_valid) begin
              pending_6 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_5_valid) begin
            pending_6 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_5_valid) begin
          pending_6 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_7 <= T_733_7;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h7 == myMaxDev) begin
            pending_7 <= GEN_2;
          end else begin
            if(io_devices_6_valid) begin
              pending_7 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_6_valid) begin
            pending_7 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_6_valid) begin
          pending_7 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_8 <= T_733_8;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h8 == myMaxDev) begin
            pending_8 <= GEN_2;
          end else begin
            if(io_devices_7_valid) begin
              pending_8 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_7_valid) begin
            pending_8 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_7_valid) begin
          pending_8 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_9 <= T_733_9;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h9 == myMaxDev) begin
            pending_9 <= GEN_2;
          end else begin
            if(io_devices_8_valid) begin
              pending_9 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_8_valid) begin
            pending_9 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_8_valid) begin
          pending_9 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_10 <= T_733_10;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'ha == myMaxDev) begin
            pending_10 <= GEN_2;
          end else begin
            if(io_devices_9_valid) begin
              pending_10 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_9_valid) begin
            pending_10 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_9_valid) begin
          pending_10 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_11 <= T_733_11;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'hb == myMaxDev) begin
            pending_11 <= GEN_2;
          end else begin
            if(io_devices_10_valid) begin
              pending_11 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_10_valid) begin
            pending_11 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_10_valid) begin
          pending_11 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_12 <= T_733_12;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'hc == myMaxDev) begin
            pending_12 <= GEN_2;
          end else begin
            if(io_devices_11_valid) begin
              pending_12 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_11_valid) begin
            pending_12 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_11_valid) begin
          pending_12 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_13 <= T_733_13;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'hd == myMaxDev) begin
            pending_13 <= GEN_2;
          end else begin
            if(io_devices_12_valid) begin
              pending_13 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_12_valid) begin
            pending_13 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_12_valid) begin
          pending_13 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_14 <= T_733_14;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'he == myMaxDev) begin
            pending_14 <= GEN_2;
          end else begin
            if(io_devices_13_valid) begin
              pending_14 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_13_valid) begin
            pending_14 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_13_valid) begin
          pending_14 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_15 <= T_733_15;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'hf == myMaxDev) begin
            pending_15 <= GEN_2;
          end else begin
            if(io_devices_14_valid) begin
              pending_15 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_14_valid) begin
            pending_15 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_14_valid) begin
          pending_15 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_16 <= T_733_16;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h10 == myMaxDev) begin
            pending_16 <= GEN_2;
          end else begin
            if(io_devices_15_valid) begin
              pending_16 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_15_valid) begin
            pending_16 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_15_valid) begin
          pending_16 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_17 <= T_733_17;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h11 == myMaxDev) begin
            pending_17 <= GEN_2;
          end else begin
            if(io_devices_16_valid) begin
              pending_17 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_16_valid) begin
            pending_17 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_16_valid) begin
          pending_17 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_18 <= T_733_18;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h12 == myMaxDev) begin
            pending_18 <= GEN_2;
          end else begin
            if(io_devices_17_valid) begin
              pending_18 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_17_valid) begin
            pending_18 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_17_valid) begin
          pending_18 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_19 <= T_733_19;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h13 == myMaxDev) begin
            pending_19 <= GEN_2;
          end else begin
            if(io_devices_18_valid) begin
              pending_19 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_18_valid) begin
            pending_19 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_18_valid) begin
          pending_19 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_20 <= T_733_20;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h14 == myMaxDev) begin
            pending_20 <= GEN_2;
          end else begin
            if(io_devices_19_valid) begin
              pending_20 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_19_valid) begin
            pending_20 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_19_valid) begin
          pending_20 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_21 <= T_733_21;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h15 == myMaxDev) begin
            pending_21 <= GEN_2;
          end else begin
            if(io_devices_20_valid) begin
              pending_21 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_20_valid) begin
            pending_21 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_20_valid) begin
          pending_21 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_22 <= T_733_22;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h16 == myMaxDev) begin
            pending_22 <= GEN_2;
          end else begin
            if(io_devices_21_valid) begin
              pending_22 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_21_valid) begin
            pending_22 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_21_valid) begin
          pending_22 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_23 <= T_733_23;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h17 == myMaxDev) begin
            pending_23 <= GEN_2;
          end else begin
            if(io_devices_22_valid) begin
              pending_23 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_22_valid) begin
            pending_23 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_22_valid) begin
          pending_23 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_24 <= T_733_24;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h18 == myMaxDev) begin
            pending_24 <= GEN_2;
          end else begin
            if(io_devices_23_valid) begin
              pending_24 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_23_valid) begin
            pending_24 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_23_valid) begin
          pending_24 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_25 <= T_733_25;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h19 == myMaxDev) begin
            pending_25 <= GEN_2;
          end else begin
            if(io_devices_24_valid) begin
              pending_25 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_24_valid) begin
            pending_25 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_24_valid) begin
          pending_25 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_26 <= T_733_26;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h1a == myMaxDev) begin
            pending_26 <= GEN_2;
          end else begin
            if(io_devices_25_valid) begin
              pending_26 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_25_valid) begin
            pending_26 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_25_valid) begin
          pending_26 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_27 <= T_733_27;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h1b == myMaxDev) begin
            pending_27 <= GEN_2;
          end else begin
            if(io_devices_26_valid) begin
              pending_27 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_26_valid) begin
            pending_27 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_26_valid) begin
          pending_27 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_28 <= T_733_28;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h1c == myMaxDev) begin
            pending_28 <= GEN_2;
          end else begin
            if(io_devices_27_valid) begin
              pending_28 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_27_valid) begin
            pending_28 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_27_valid) begin
          pending_28 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_29 <= T_733_29;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h1d == myMaxDev) begin
            pending_29 <= GEN_2;
          end else begin
            if(io_devices_28_valid) begin
              pending_29 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_28_valid) begin
            pending_29 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_28_valid) begin
          pending_29 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_30 <= T_733_30;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h1e == myMaxDev) begin
            pending_30 <= GEN_2;
          end else begin
            if(io_devices_29_valid) begin
              pending_30 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_29_valid) begin
            pending_30 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_29_valid) begin
          pending_30 <= 1'h1;
        end
      end
    end
    if(reset) begin
      pending_31 <= T_733_31;
    end else begin
      if(T_1406) begin
        if(T_1415) begin
          if(5'h1f == myMaxDev) begin
            pending_31 <= GEN_2;
          end else begin
            if(io_devices_30_valid) begin
              pending_31 <= 1'h1;
            end
          end
        end else begin
          if(io_devices_30_valid) begin
            pending_31 <= 1'h1;
          end
        end
      end else begin
        if(io_devices_30_valid) begin
          pending_31 <= 1'h1;
        end
      end
    end
    if(1'h0) begin
    end else begin
      enables_0_0 <= 1'h0;
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_1 <= GEN_38;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_2 <= GEN_39;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_3 <= GEN_40;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_4 <= GEN_41;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_5 <= GEN_42;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_6 <= GEN_43;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_7 <= GEN_44;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_8 <= GEN_45;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_9 <= GEN_46;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_10 <= GEN_47;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_11 <= GEN_48;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_12 <= GEN_49;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_13 <= GEN_50;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_14 <= GEN_51;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_15 <= GEN_52;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_16 <= GEN_53;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_17 <= GEN_54;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_18 <= GEN_55;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_19 <= GEN_56;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_20 <= GEN_57;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_21 <= GEN_58;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_22 <= GEN_59;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_23 <= GEN_60;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_24 <= GEN_61;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_25 <= GEN_62;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_26 <= GEN_63;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_27 <= GEN_64;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_28 <= GEN_65;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_29 <= GEN_66;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_30 <= GEN_67;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1462) begin
        if(write) begin
          enables_0_31 <= GEN_68;
        end
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1176) begin
        T_1182 <= {{1'd0}, T_1069};
      end else begin
        T_1182 <= T_1180;
      end
    end
    if(1'h0) begin
    end else begin
      if(T_1176) begin
        if(T_1064) begin
          if(T_1008) begin
            if(T_980) begin
              if(T_966) begin
                T_1183 <= 2'h2;
              end else begin
                T_1183 <= T_901;
              end
            end else begin
              if(T_974) begin
                T_1183 <= T_903;
              end else begin
                T_1183 <= T_905;
              end
            end
          end else begin
            if(T_1002) begin
              if(T_988) begin
                T_1183 <= T_907;
              end else begin
                T_1183 <= T_909;
              end
            end else begin
              if(T_996) begin
                T_1183 <= T_911;
              end else begin
                T_1183 <= T_913;
              end
            end
          end
        end else begin
          if(T_1058) begin
            if(T_1030) begin
              if(T_1016) begin
                T_1183 <= T_915;
              end else begin
                T_1183 <= T_917;
              end
            end else begin
              if(T_1024) begin
                T_1183 <= T_919;
              end else begin
                T_1183 <= T_921;
              end
            end
          end else begin
            if(T_1052) begin
              if(T_1038) begin
                T_1183 <= T_923;
              end else begin
                T_1183 <= T_925;
              end
            end else begin
              if(T_1046) begin
                T_1183 <= T_927;
              end else begin
                T_1183 <= T_929;
              end
            end
          end
        end
      end else begin
        if(T_1170) begin
          if(T_1114) begin
            if(T_1086) begin
              if(T_1072) begin
                T_1183 <= T_931;
              end else begin
                T_1183 <= T_933;
              end
            end else begin
              if(T_1080) begin
                T_1183 <= T_935;
              end else begin
                T_1183 <= T_937;
              end
            end
          end else begin
            if(T_1108) begin
              if(T_1094) begin
                T_1183 <= T_939;
              end else begin
                T_1183 <= T_941;
              end
            end else begin
              if(T_1102) begin
                T_1183 <= T_943;
              end else begin
                T_1183 <= T_945;
              end
            end
          end
        end else begin
          if(T_1164) begin
            if(T_1136) begin
              if(T_1122) begin
                T_1183 <= T_947;
              end else begin
                T_1183 <= T_949;
              end
            end else begin
              if(T_1130) begin
                T_1183 <= T_951;
              end else begin
                T_1183 <= T_953;
              end
            end
          end else begin
            if(T_1158) begin
              if(T_1144) begin
                T_1183 <= T_955;
              end else begin
                T_1183 <= T_957;
              end
            end else begin
              if(T_1152) begin
                T_1183 <= T_959;
              end else begin
                T_1183 <= T_961;
              end
            end
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (T_1225) begin
          $fwrite(32'h80000002,"Assertion failed: unsupported PLIC operation\n    at Plic.scala:108 assert(!acq.fire() || read || write, ---unsupported PLIC operation---)\n");
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (T_1225) begin
          $fatal;
        end
    `ifdef STOP_COND
      end
    `endif
    `endif
  end
endmodule
